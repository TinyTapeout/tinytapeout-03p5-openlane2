module tt_mux (k_one,
    k_zero,
    addr,
    spine_iw,
    spine_ow,
    um_ena,
    um_iw,
    um_k_zero,
    um_ow);
 output k_one;
 output k_zero;
 input [4:0] addr;
 input [30:0] spine_iw;
 output [25:0] spine_ow;
 output [15:0] um_ena;
 output [287:0] um_iw;
 output [15:0] um_k_zero;
 input [383:0] um_ow;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire \col[0].genblk1.mux4_I[0].x ;
 wire \col[0].genblk1.mux4_I[10].x ;
 wire \col[0].genblk1.mux4_I[11].x ;
 wire \col[0].genblk1.mux4_I[12].x ;
 wire \col[0].genblk1.mux4_I[13].x ;
 wire \col[0].genblk1.mux4_I[14].x ;
 wire \col[0].genblk1.mux4_I[15].x ;
 wire \col[0].genblk1.mux4_I[16].x ;
 wire \col[0].genblk1.mux4_I[17].x ;
 wire \col[0].genblk1.mux4_I[18].x ;
 wire \col[0].genblk1.mux4_I[19].x ;
 wire \col[0].genblk1.mux4_I[1].x ;
 wire \col[0].genblk1.mux4_I[20].x ;
 wire \col[0].genblk1.mux4_I[21].x ;
 wire \col[0].genblk1.mux4_I[22].x ;
 wire \col[0].genblk1.mux4_I[23].x ;
 wire \col[0].genblk1.mux4_I[2].x ;
 wire \col[0].genblk1.mux4_I[3].x ;
 wire \col[0].genblk1.mux4_I[4].x ;
 wire \col[0].genblk1.mux4_I[5].x ;
 wire \col[0].genblk1.mux4_I[6].x ;
 wire \col[0].genblk1.mux4_I[7].x ;
 wire \col[0].genblk1.mux4_I[8].x ;
 wire \col[0].genblk1.mux4_I[9].x ;
 wire \col[0].genblk1.tbuf_row_ena_I.t ;
 wire \col[0].genblk1.tbuf_row_ena_I.tx ;
 wire \col[0].genblk1.tbuf_spine_ow_I[0].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[10].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[11].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[12].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[13].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[14].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[15].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[16].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[17].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[18].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[19].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[1].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[20].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[21].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[22].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[23].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[2].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[3].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[4].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[5].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[6].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[7].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[8].z ;
 wire \col[0].genblk1.tbuf_spine_ow_I[9].z ;
 wire \col[0].tie_bot_I.hi ;
 wire \col[0].tie_bot_I.lo ;
 wire \col[0].tie_top_I.hi ;
 wire \col[0].tie_top_I.lo ;
 wire \col[0].zbuf_bot_ena_I.e ;
 wire \col[0].zbuf_bot_ena_I.z ;
 wire \col[0].zbuf_bot_iw_I[0].a ;
 wire \col[0].zbuf_bot_iw_I[0].z ;
 wire \col[0].zbuf_bot_iw_I[10].a ;
 wire \col[0].zbuf_bot_iw_I[10].z ;
 wire \col[0].zbuf_bot_iw_I[11].a ;
 wire \col[0].zbuf_bot_iw_I[11].z ;
 wire \col[0].zbuf_bot_iw_I[12].a ;
 wire \col[0].zbuf_bot_iw_I[12].z ;
 wire \col[0].zbuf_bot_iw_I[13].a ;
 wire \col[0].zbuf_bot_iw_I[13].z ;
 wire \col[0].zbuf_bot_iw_I[14].a ;
 wire \col[0].zbuf_bot_iw_I[14].z ;
 wire \col[0].zbuf_bot_iw_I[15].a ;
 wire \col[0].zbuf_bot_iw_I[15].z ;
 wire \col[0].zbuf_bot_iw_I[16].a ;
 wire \col[0].zbuf_bot_iw_I[16].z ;
 wire \col[0].zbuf_bot_iw_I[17].a ;
 wire \col[0].zbuf_bot_iw_I[17].z ;
 wire \col[0].zbuf_bot_iw_I[1].a ;
 wire \col[0].zbuf_bot_iw_I[1].z ;
 wire \col[0].zbuf_bot_iw_I[2].a ;
 wire \col[0].zbuf_bot_iw_I[2].z ;
 wire \col[0].zbuf_bot_iw_I[3].a ;
 wire \col[0].zbuf_bot_iw_I[3].z ;
 wire \col[0].zbuf_bot_iw_I[4].a ;
 wire \col[0].zbuf_bot_iw_I[4].z ;
 wire \col[0].zbuf_bot_iw_I[5].a ;
 wire \col[0].zbuf_bot_iw_I[5].z ;
 wire \col[0].zbuf_bot_iw_I[6].a ;
 wire \col[0].zbuf_bot_iw_I[6].z ;
 wire \col[0].zbuf_bot_iw_I[7].a ;
 wire \col[0].zbuf_bot_iw_I[7].z ;
 wire \col[0].zbuf_bot_iw_I[8].a ;
 wire \col[0].zbuf_bot_iw_I[8].z ;
 wire \col[0].zbuf_bot_iw_I[9].a ;
 wire \col[0].zbuf_bot_iw_I[9].z ;
 wire \col[0].zbuf_top_ena_I.e ;
 wire \col[0].zbuf_top_ena_I.z ;
 wire \col[0].zbuf_top_iw_I[0].z ;
 wire \col[0].zbuf_top_iw_I[10].z ;
 wire \col[0].zbuf_top_iw_I[11].z ;
 wire \col[0].zbuf_top_iw_I[12].z ;
 wire \col[0].zbuf_top_iw_I[13].z ;
 wire \col[0].zbuf_top_iw_I[14].z ;
 wire \col[0].zbuf_top_iw_I[15].z ;
 wire \col[0].zbuf_top_iw_I[16].z ;
 wire \col[0].zbuf_top_iw_I[17].z ;
 wire \col[0].zbuf_top_iw_I[1].z ;
 wire \col[0].zbuf_top_iw_I[2].z ;
 wire \col[0].zbuf_top_iw_I[3].z ;
 wire \col[0].zbuf_top_iw_I[4].z ;
 wire \col[0].zbuf_top_iw_I[5].z ;
 wire \col[0].zbuf_top_iw_I[6].z ;
 wire \col[0].zbuf_top_iw_I[7].z ;
 wire \col[0].zbuf_top_iw_I[8].z ;
 wire \col[0].zbuf_top_iw_I[9].z ;
 wire \col[1].tie_bot_I.hi ;
 wire \col[1].tie_bot_I.lo ;
 wire \col[1].tie_top_I.hi ;
 wire \col[1].tie_top_I.lo ;
 wire \col[1].zbuf_bot_ena_I.e ;
 wire \col[1].zbuf_bot_ena_I.z ;
 wire \col[1].zbuf_bot_iw_I[0].z ;
 wire \col[1].zbuf_bot_iw_I[10].z ;
 wire \col[1].zbuf_bot_iw_I[11].z ;
 wire \col[1].zbuf_bot_iw_I[12].z ;
 wire \col[1].zbuf_bot_iw_I[13].z ;
 wire \col[1].zbuf_bot_iw_I[14].z ;
 wire \col[1].zbuf_bot_iw_I[15].z ;
 wire \col[1].zbuf_bot_iw_I[16].z ;
 wire \col[1].zbuf_bot_iw_I[17].z ;
 wire \col[1].zbuf_bot_iw_I[1].z ;
 wire \col[1].zbuf_bot_iw_I[2].z ;
 wire \col[1].zbuf_bot_iw_I[3].z ;
 wire \col[1].zbuf_bot_iw_I[4].z ;
 wire \col[1].zbuf_bot_iw_I[5].z ;
 wire \col[1].zbuf_bot_iw_I[6].z ;
 wire \col[1].zbuf_bot_iw_I[7].z ;
 wire \col[1].zbuf_bot_iw_I[8].z ;
 wire \col[1].zbuf_bot_iw_I[9].z ;
 wire \col[1].zbuf_top_ena_I.e ;
 wire \col[1].zbuf_top_ena_I.z ;
 wire \col[1].zbuf_top_iw_I[0].z ;
 wire \col[1].zbuf_top_iw_I[10].z ;
 wire \col[1].zbuf_top_iw_I[11].z ;
 wire \col[1].zbuf_top_iw_I[12].z ;
 wire \col[1].zbuf_top_iw_I[13].z ;
 wire \col[1].zbuf_top_iw_I[14].z ;
 wire \col[1].zbuf_top_iw_I[15].z ;
 wire \col[1].zbuf_top_iw_I[16].z ;
 wire \col[1].zbuf_top_iw_I[17].z ;
 wire \col[1].zbuf_top_iw_I[1].z ;
 wire \col[1].zbuf_top_iw_I[2].z ;
 wire \col[1].zbuf_top_iw_I[3].z ;
 wire \col[1].zbuf_top_iw_I[4].z ;
 wire \col[1].zbuf_top_iw_I[5].z ;
 wire \col[1].zbuf_top_iw_I[6].z ;
 wire \col[1].zbuf_top_iw_I[7].z ;
 wire \col[1].zbuf_top_iw_I[8].z ;
 wire \col[1].zbuf_top_iw_I[9].z ;
 wire \col[2].genblk1.mux4_I[0].x ;
 wire \col[2].genblk1.mux4_I[10].x ;
 wire \col[2].genblk1.mux4_I[11].x ;
 wire \col[2].genblk1.mux4_I[12].x ;
 wire \col[2].genblk1.mux4_I[13].x ;
 wire \col[2].genblk1.mux4_I[14].x ;
 wire \col[2].genblk1.mux4_I[15].x ;
 wire \col[2].genblk1.mux4_I[16].x ;
 wire \col[2].genblk1.mux4_I[17].x ;
 wire \col[2].genblk1.mux4_I[18].x ;
 wire \col[2].genblk1.mux4_I[19].x ;
 wire \col[2].genblk1.mux4_I[1].x ;
 wire \col[2].genblk1.mux4_I[20].x ;
 wire \col[2].genblk1.mux4_I[21].x ;
 wire \col[2].genblk1.mux4_I[22].x ;
 wire \col[2].genblk1.mux4_I[23].x ;
 wire \col[2].genblk1.mux4_I[2].x ;
 wire \col[2].genblk1.mux4_I[3].x ;
 wire \col[2].genblk1.mux4_I[4].x ;
 wire \col[2].genblk1.mux4_I[5].x ;
 wire \col[2].genblk1.mux4_I[6].x ;
 wire \col[2].genblk1.mux4_I[7].x ;
 wire \col[2].genblk1.mux4_I[8].x ;
 wire \col[2].genblk1.mux4_I[9].x ;
 wire \col[2].genblk1.tbuf_row_ena_I.t ;
 wire \col[2].genblk1.tbuf_row_ena_I.tx ;
 wire \col[2].tie_bot_I.hi ;
 wire \col[2].tie_bot_I.lo ;
 wire \col[2].tie_top_I.hi ;
 wire \col[2].tie_top_I.lo ;
 wire \col[2].zbuf_bot_ena_I.e ;
 wire \col[2].zbuf_bot_ena_I.z ;
 wire \col[2].zbuf_bot_iw_I[0].z ;
 wire \col[2].zbuf_bot_iw_I[10].z ;
 wire \col[2].zbuf_bot_iw_I[11].z ;
 wire \col[2].zbuf_bot_iw_I[12].z ;
 wire \col[2].zbuf_bot_iw_I[13].z ;
 wire \col[2].zbuf_bot_iw_I[14].z ;
 wire \col[2].zbuf_bot_iw_I[15].z ;
 wire \col[2].zbuf_bot_iw_I[16].z ;
 wire \col[2].zbuf_bot_iw_I[17].z ;
 wire \col[2].zbuf_bot_iw_I[1].z ;
 wire \col[2].zbuf_bot_iw_I[2].z ;
 wire \col[2].zbuf_bot_iw_I[3].z ;
 wire \col[2].zbuf_bot_iw_I[4].z ;
 wire \col[2].zbuf_bot_iw_I[5].z ;
 wire \col[2].zbuf_bot_iw_I[6].z ;
 wire \col[2].zbuf_bot_iw_I[7].z ;
 wire \col[2].zbuf_bot_iw_I[8].z ;
 wire \col[2].zbuf_bot_iw_I[9].z ;
 wire \col[2].zbuf_top_ena_I.e ;
 wire \col[2].zbuf_top_ena_I.z ;
 wire \col[2].zbuf_top_iw_I[0].z ;
 wire \col[2].zbuf_top_iw_I[10].z ;
 wire \col[2].zbuf_top_iw_I[11].z ;
 wire \col[2].zbuf_top_iw_I[12].z ;
 wire \col[2].zbuf_top_iw_I[13].z ;
 wire \col[2].zbuf_top_iw_I[14].z ;
 wire \col[2].zbuf_top_iw_I[15].z ;
 wire \col[2].zbuf_top_iw_I[16].z ;
 wire \col[2].zbuf_top_iw_I[17].z ;
 wire \col[2].zbuf_top_iw_I[1].z ;
 wire \col[2].zbuf_top_iw_I[2].z ;
 wire \col[2].zbuf_top_iw_I[3].z ;
 wire \col[2].zbuf_top_iw_I[4].z ;
 wire \col[2].zbuf_top_iw_I[5].z ;
 wire \col[2].zbuf_top_iw_I[6].z ;
 wire \col[2].zbuf_top_iw_I[7].z ;
 wire \col[2].zbuf_top_iw_I[8].z ;
 wire \col[2].zbuf_top_iw_I[9].z ;
 wire \col[3].tie_bot_I.hi ;
 wire \col[3].tie_bot_I.lo ;
 wire \col[3].tie_top_I.hi ;
 wire \col[3].tie_top_I.lo ;
 wire \col[3].zbuf_bot_ena_I.e ;
 wire \col[3].zbuf_bot_ena_I.z ;
 wire \col[3].zbuf_bot_iw_I[0].z ;
 wire \col[3].zbuf_bot_iw_I[10].z ;
 wire \col[3].zbuf_bot_iw_I[11].z ;
 wire \col[3].zbuf_bot_iw_I[12].z ;
 wire \col[3].zbuf_bot_iw_I[13].z ;
 wire \col[3].zbuf_bot_iw_I[14].z ;
 wire \col[3].zbuf_bot_iw_I[15].z ;
 wire \col[3].zbuf_bot_iw_I[16].z ;
 wire \col[3].zbuf_bot_iw_I[17].z ;
 wire \col[3].zbuf_bot_iw_I[1].z ;
 wire \col[3].zbuf_bot_iw_I[2].z ;
 wire \col[3].zbuf_bot_iw_I[3].z ;
 wire \col[3].zbuf_bot_iw_I[4].z ;
 wire \col[3].zbuf_bot_iw_I[5].z ;
 wire \col[3].zbuf_bot_iw_I[6].z ;
 wire \col[3].zbuf_bot_iw_I[7].z ;
 wire \col[3].zbuf_bot_iw_I[8].z ;
 wire \col[3].zbuf_bot_iw_I[9].z ;
 wire \col[3].zbuf_top_ena_I.e ;
 wire \col[3].zbuf_top_ena_I.z ;
 wire \col[3].zbuf_top_iw_I[0].z ;
 wire \col[3].zbuf_top_iw_I[10].z ;
 wire \col[3].zbuf_top_iw_I[11].z ;
 wire \col[3].zbuf_top_iw_I[12].z ;
 wire \col[3].zbuf_top_iw_I[13].z ;
 wire \col[3].zbuf_top_iw_I[14].z ;
 wire \col[3].zbuf_top_iw_I[15].z ;
 wire \col[3].zbuf_top_iw_I[16].z ;
 wire \col[3].zbuf_top_iw_I[17].z ;
 wire \col[3].zbuf_top_iw_I[1].z ;
 wire \col[3].zbuf_top_iw_I[2].z ;
 wire \col[3].zbuf_top_iw_I[3].z ;
 wire \col[3].zbuf_top_iw_I[4].z ;
 wire \col[3].zbuf_top_iw_I[5].z ;
 wire \col[3].zbuf_top_iw_I[6].z ;
 wire \col[3].zbuf_top_iw_I[7].z ;
 wire \col[3].zbuf_top_iw_I[8].z ;
 wire \col[3].zbuf_top_iw_I[9].z ;
 wire \col[4].genblk1.mux4_I[0].x ;
 wire \col[4].genblk1.mux4_I[10].x ;
 wire \col[4].genblk1.mux4_I[11].x ;
 wire \col[4].genblk1.mux4_I[12].x ;
 wire \col[4].genblk1.mux4_I[13].x ;
 wire \col[4].genblk1.mux4_I[14].x ;
 wire \col[4].genblk1.mux4_I[15].x ;
 wire \col[4].genblk1.mux4_I[16].x ;
 wire \col[4].genblk1.mux4_I[17].x ;
 wire \col[4].genblk1.mux4_I[18].x ;
 wire \col[4].genblk1.mux4_I[19].x ;
 wire \col[4].genblk1.mux4_I[1].x ;
 wire \col[4].genblk1.mux4_I[20].x ;
 wire \col[4].genblk1.mux4_I[21].x ;
 wire \col[4].genblk1.mux4_I[22].x ;
 wire \col[4].genblk1.mux4_I[23].x ;
 wire \col[4].genblk1.mux4_I[2].x ;
 wire \col[4].genblk1.mux4_I[3].x ;
 wire \col[4].genblk1.mux4_I[4].x ;
 wire \col[4].genblk1.mux4_I[5].x ;
 wire \col[4].genblk1.mux4_I[6].x ;
 wire \col[4].genblk1.mux4_I[7].x ;
 wire \col[4].genblk1.mux4_I[8].x ;
 wire \col[4].genblk1.mux4_I[9].x ;
 wire \col[4].genblk1.tbuf_row_ena_I.t ;
 wire \col[4].genblk1.tbuf_row_ena_I.tx ;
 wire \col[4].tie_bot_I.hi ;
 wire \col[4].tie_bot_I.lo ;
 wire \col[4].tie_top_I.hi ;
 wire \col[4].tie_top_I.lo ;
 wire \col[4].zbuf_bot_ena_I.e ;
 wire \col[4].zbuf_bot_ena_I.z ;
 wire \col[4].zbuf_bot_iw_I[0].z ;
 wire \col[4].zbuf_bot_iw_I[10].z ;
 wire \col[4].zbuf_bot_iw_I[11].z ;
 wire \col[4].zbuf_bot_iw_I[12].z ;
 wire \col[4].zbuf_bot_iw_I[13].z ;
 wire \col[4].zbuf_bot_iw_I[14].z ;
 wire \col[4].zbuf_bot_iw_I[15].z ;
 wire \col[4].zbuf_bot_iw_I[16].z ;
 wire \col[4].zbuf_bot_iw_I[17].z ;
 wire \col[4].zbuf_bot_iw_I[1].z ;
 wire \col[4].zbuf_bot_iw_I[2].z ;
 wire \col[4].zbuf_bot_iw_I[3].z ;
 wire \col[4].zbuf_bot_iw_I[4].z ;
 wire \col[4].zbuf_bot_iw_I[5].z ;
 wire \col[4].zbuf_bot_iw_I[6].z ;
 wire \col[4].zbuf_bot_iw_I[7].z ;
 wire \col[4].zbuf_bot_iw_I[8].z ;
 wire \col[4].zbuf_bot_iw_I[9].z ;
 wire \col[4].zbuf_top_ena_I.e ;
 wire \col[4].zbuf_top_ena_I.z ;
 wire \col[4].zbuf_top_iw_I[0].z ;
 wire \col[4].zbuf_top_iw_I[10].z ;
 wire \col[4].zbuf_top_iw_I[11].z ;
 wire \col[4].zbuf_top_iw_I[12].z ;
 wire \col[4].zbuf_top_iw_I[13].z ;
 wire \col[4].zbuf_top_iw_I[14].z ;
 wire \col[4].zbuf_top_iw_I[15].z ;
 wire \col[4].zbuf_top_iw_I[16].z ;
 wire \col[4].zbuf_top_iw_I[17].z ;
 wire \col[4].zbuf_top_iw_I[1].z ;
 wire \col[4].zbuf_top_iw_I[2].z ;
 wire \col[4].zbuf_top_iw_I[3].z ;
 wire \col[4].zbuf_top_iw_I[4].z ;
 wire \col[4].zbuf_top_iw_I[5].z ;
 wire \col[4].zbuf_top_iw_I[6].z ;
 wire \col[4].zbuf_top_iw_I[7].z ;
 wire \col[4].zbuf_top_iw_I[8].z ;
 wire \col[4].zbuf_top_iw_I[9].z ;
 wire \col[5].tie_bot_I.hi ;
 wire \col[5].tie_bot_I.lo ;
 wire \col[5].tie_top_I.hi ;
 wire \col[5].tie_top_I.lo ;
 wire \col[5].zbuf_bot_ena_I.e ;
 wire \col[5].zbuf_bot_ena_I.z ;
 wire \col[5].zbuf_bot_iw_I[0].z ;
 wire \col[5].zbuf_bot_iw_I[10].z ;
 wire \col[5].zbuf_bot_iw_I[11].z ;
 wire \col[5].zbuf_bot_iw_I[12].z ;
 wire \col[5].zbuf_bot_iw_I[13].z ;
 wire \col[5].zbuf_bot_iw_I[14].z ;
 wire \col[5].zbuf_bot_iw_I[15].z ;
 wire \col[5].zbuf_bot_iw_I[16].z ;
 wire \col[5].zbuf_bot_iw_I[17].z ;
 wire \col[5].zbuf_bot_iw_I[1].z ;
 wire \col[5].zbuf_bot_iw_I[2].z ;
 wire \col[5].zbuf_bot_iw_I[3].z ;
 wire \col[5].zbuf_bot_iw_I[4].z ;
 wire \col[5].zbuf_bot_iw_I[5].z ;
 wire \col[5].zbuf_bot_iw_I[6].z ;
 wire \col[5].zbuf_bot_iw_I[7].z ;
 wire \col[5].zbuf_bot_iw_I[8].z ;
 wire \col[5].zbuf_bot_iw_I[9].z ;
 wire \col[5].zbuf_top_ena_I.e ;
 wire \col[5].zbuf_top_ena_I.z ;
 wire \col[5].zbuf_top_iw_I[0].z ;
 wire \col[5].zbuf_top_iw_I[10].z ;
 wire \col[5].zbuf_top_iw_I[11].z ;
 wire \col[5].zbuf_top_iw_I[12].z ;
 wire \col[5].zbuf_top_iw_I[13].z ;
 wire \col[5].zbuf_top_iw_I[14].z ;
 wire \col[5].zbuf_top_iw_I[15].z ;
 wire \col[5].zbuf_top_iw_I[16].z ;
 wire \col[5].zbuf_top_iw_I[17].z ;
 wire \col[5].zbuf_top_iw_I[1].z ;
 wire \col[5].zbuf_top_iw_I[2].z ;
 wire \col[5].zbuf_top_iw_I[3].z ;
 wire \col[5].zbuf_top_iw_I[4].z ;
 wire \col[5].zbuf_top_iw_I[5].z ;
 wire \col[5].zbuf_top_iw_I[6].z ;
 wire \col[5].zbuf_top_iw_I[7].z ;
 wire \col[5].zbuf_top_iw_I[8].z ;
 wire \col[5].zbuf_top_iw_I[9].z ;
 wire \col[6].genblk1.mux4_I[0].x ;
 wire \col[6].genblk1.mux4_I[10].x ;
 wire \col[6].genblk1.mux4_I[11].x ;
 wire \col[6].genblk1.mux4_I[12].x ;
 wire \col[6].genblk1.mux4_I[13].x ;
 wire \col[6].genblk1.mux4_I[14].x ;
 wire \col[6].genblk1.mux4_I[15].x ;
 wire \col[6].genblk1.mux4_I[16].x ;
 wire \col[6].genblk1.mux4_I[17].x ;
 wire \col[6].genblk1.mux4_I[18].x ;
 wire \col[6].genblk1.mux4_I[19].x ;
 wire \col[6].genblk1.mux4_I[1].x ;
 wire \col[6].genblk1.mux4_I[20].x ;
 wire \col[6].genblk1.mux4_I[21].x ;
 wire \col[6].genblk1.mux4_I[22].x ;
 wire \col[6].genblk1.mux4_I[23].x ;
 wire \col[6].genblk1.mux4_I[2].x ;
 wire \col[6].genblk1.mux4_I[3].x ;
 wire \col[6].genblk1.mux4_I[4].x ;
 wire \col[6].genblk1.mux4_I[5].x ;
 wire \col[6].genblk1.mux4_I[6].x ;
 wire \col[6].genblk1.mux4_I[7].x ;
 wire \col[6].genblk1.mux4_I[8].x ;
 wire \col[6].genblk1.mux4_I[9].x ;
 wire \col[6].genblk1.tbuf_row_ena_I.t ;
 wire \col[6].genblk1.tbuf_row_ena_I.tx ;
 wire \col[6].tie_bot_I.hi ;
 wire \col[6].tie_bot_I.lo ;
 wire \col[6].tie_top_I.hi ;
 wire \col[6].tie_top_I.lo ;
 wire \col[6].zbuf_bot_ena_I.e ;
 wire \col[6].zbuf_bot_ena_I.z ;
 wire \col[6].zbuf_bot_iw_I[0].z ;
 wire \col[6].zbuf_bot_iw_I[10].z ;
 wire \col[6].zbuf_bot_iw_I[11].z ;
 wire \col[6].zbuf_bot_iw_I[12].z ;
 wire \col[6].zbuf_bot_iw_I[13].z ;
 wire \col[6].zbuf_bot_iw_I[14].z ;
 wire \col[6].zbuf_bot_iw_I[15].z ;
 wire \col[6].zbuf_bot_iw_I[16].z ;
 wire \col[6].zbuf_bot_iw_I[17].z ;
 wire \col[6].zbuf_bot_iw_I[1].z ;
 wire \col[6].zbuf_bot_iw_I[2].z ;
 wire \col[6].zbuf_bot_iw_I[3].z ;
 wire \col[6].zbuf_bot_iw_I[4].z ;
 wire \col[6].zbuf_bot_iw_I[5].z ;
 wire \col[6].zbuf_bot_iw_I[6].z ;
 wire \col[6].zbuf_bot_iw_I[7].z ;
 wire \col[6].zbuf_bot_iw_I[8].z ;
 wire \col[6].zbuf_bot_iw_I[9].z ;
 wire \col[6].zbuf_top_ena_I.e ;
 wire \col[6].zbuf_top_ena_I.z ;
 wire \col[6].zbuf_top_iw_I[0].z ;
 wire \col[6].zbuf_top_iw_I[10].z ;
 wire \col[6].zbuf_top_iw_I[11].z ;
 wire \col[6].zbuf_top_iw_I[12].z ;
 wire \col[6].zbuf_top_iw_I[13].z ;
 wire \col[6].zbuf_top_iw_I[14].z ;
 wire \col[6].zbuf_top_iw_I[15].z ;
 wire \col[6].zbuf_top_iw_I[16].z ;
 wire \col[6].zbuf_top_iw_I[17].z ;
 wire \col[6].zbuf_top_iw_I[1].z ;
 wire \col[6].zbuf_top_iw_I[2].z ;
 wire \col[6].zbuf_top_iw_I[3].z ;
 wire \col[6].zbuf_top_iw_I[4].z ;
 wire \col[6].zbuf_top_iw_I[5].z ;
 wire \col[6].zbuf_top_iw_I[6].z ;
 wire \col[6].zbuf_top_iw_I[7].z ;
 wire \col[6].zbuf_top_iw_I[8].z ;
 wire \col[6].zbuf_top_iw_I[9].z ;
 wire \col[7].tie_bot_I.hi ;
 wire \col[7].tie_bot_I.lo ;
 wire \col[7].tie_top_I.hi ;
 wire \col[7].tie_top_I.lo ;
 wire \col[7].zbuf_bot_ena_I.e ;
 wire \col[7].zbuf_bot_ena_I.z ;
 wire \col[7].zbuf_bot_iw_I[0].z ;
 wire \col[7].zbuf_bot_iw_I[10].z ;
 wire \col[7].zbuf_bot_iw_I[11].z ;
 wire \col[7].zbuf_bot_iw_I[12].z ;
 wire \col[7].zbuf_bot_iw_I[13].z ;
 wire \col[7].zbuf_bot_iw_I[14].z ;
 wire \col[7].zbuf_bot_iw_I[15].z ;
 wire \col[7].zbuf_bot_iw_I[16].z ;
 wire \col[7].zbuf_bot_iw_I[17].z ;
 wire \col[7].zbuf_bot_iw_I[1].z ;
 wire \col[7].zbuf_bot_iw_I[2].z ;
 wire \col[7].zbuf_bot_iw_I[3].z ;
 wire \col[7].zbuf_bot_iw_I[4].z ;
 wire \col[7].zbuf_bot_iw_I[5].z ;
 wire \col[7].zbuf_bot_iw_I[6].z ;
 wire \col[7].zbuf_bot_iw_I[7].z ;
 wire \col[7].zbuf_bot_iw_I[8].z ;
 wire \col[7].zbuf_bot_iw_I[9].z ;
 wire \col[7].zbuf_top_ena_I.e ;
 wire \col[7].zbuf_top_ena_I.z ;
 wire \col[7].zbuf_top_iw_I[0].z ;
 wire \col[7].zbuf_top_iw_I[10].z ;
 wire \col[7].zbuf_top_iw_I[11].z ;
 wire \col[7].zbuf_top_iw_I[12].z ;
 wire \col[7].zbuf_top_iw_I[13].z ;
 wire \col[7].zbuf_top_iw_I[14].z ;
 wire \col[7].zbuf_top_iw_I[15].z ;
 wire \col[7].zbuf_top_iw_I[16].z ;
 wire \col[7].zbuf_top_iw_I[17].z ;
 wire \col[7].zbuf_top_iw_I[1].z ;
 wire \col[7].zbuf_top_iw_I[2].z ;
 wire \col[7].zbuf_top_iw_I[3].z ;
 wire \col[7].zbuf_top_iw_I[4].z ;
 wire \col[7].zbuf_top_iw_I[5].z ;
 wire \col[7].zbuf_top_iw_I[6].z ;
 wire \col[7].zbuf_top_iw_I[7].z ;
 wire \col[7].zbuf_top_iw_I[8].z ;
 wire \col[7].zbuf_top_iw_I[9].z ;
 wire one_;
 wire \tbuf_row_ena_I.t ;
 wire \tbuf_row_ena_I.tx ;
 wire \tbuf_spine_ow_I[0].z ;
 wire \tbuf_spine_ow_I[10].z ;
 wire \tbuf_spine_ow_I[11].z ;
 wire \tbuf_spine_ow_I[12].z ;
 wire \tbuf_spine_ow_I[13].z ;
 wire \tbuf_spine_ow_I[14].z ;
 wire \tbuf_spine_ow_I[15].z ;
 wire \tbuf_spine_ow_I[16].z ;
 wire \tbuf_spine_ow_I[17].z ;
 wire \tbuf_spine_ow_I[18].z ;
 wire \tbuf_spine_ow_I[19].z ;
 wire \tbuf_spine_ow_I[1].z ;
 wire \tbuf_spine_ow_I[20].z ;
 wire \tbuf_spine_ow_I[21].z ;
 wire \tbuf_spine_ow_I[22].z ;
 wire \tbuf_spine_ow_I[23].z ;
 wire \tbuf_spine_ow_I[2].z ;
 wire \tbuf_spine_ow_I[3].z ;
 wire \tbuf_spine_ow_I[4].z ;
 wire \tbuf_spine_ow_I[5].z ;
 wire \tbuf_spine_ow_I[6].z ;
 wire \tbuf_spine_ow_I[7].z ;
 wire \tbuf_spine_ow_I[8].z ;
 wire \tbuf_spine_ow_I[9].z ;
 wire \tie_spine_guard_I[0].hi ;
 wire \tie_spine_guard_I[0].lo ;
 wire \tie_spine_guard_I[1].hi ;
 wire \tie_spine_guard_I[1].lo ;
 wire \zbuf_bus_ena_I.genblk1.l ;
 wire \zbuf_bus_ena_I.z ;
 wire \zbuf_bus_iw_I[0].genblk1.l ;
 wire \zbuf_bus_iw_I[10].genblk1.l ;
 wire \zbuf_bus_iw_I[11].genblk1.l ;
 wire \zbuf_bus_iw_I[12].genblk1.l ;
 wire \zbuf_bus_iw_I[13].genblk1.l ;
 wire \zbuf_bus_iw_I[14].genblk1.l ;
 wire \zbuf_bus_iw_I[15].genblk1.l ;
 wire \zbuf_bus_iw_I[16].genblk1.l ;
 wire \zbuf_bus_iw_I[17].genblk1.l ;
 wire \zbuf_bus_iw_I[1].genblk1.l ;
 wire \zbuf_bus_iw_I[2].genblk1.l ;
 wire \zbuf_bus_iw_I[3].genblk1.l ;
 wire \zbuf_bus_iw_I[4].genblk1.l ;
 wire \zbuf_bus_iw_I[5].genblk1.l ;
 wire \zbuf_bus_iw_I[6].genblk1.l ;
 wire \zbuf_bus_iw_I[7].genblk1.l ;
 wire \zbuf_bus_iw_I[8].genblk1.l ;
 wire \zbuf_bus_iw_I[9].genblk1.l ;
 wire \zbuf_bus_sel_I[0].genblk1.l ;
 wire \zbuf_bus_sel_I[0].z ;
 wire \zbuf_bus_sel_I[1].genblk1.l ;
 wire \zbuf_bus_sel_I[1].z ;
 wire \zbuf_bus_sel_I[2].genblk1.l ;
 wire \zbuf_bus_sel_I[2].z ;
 wire \zbuf_bus_sel_I[3].genblk1.l ;
 wire \zbuf_bus_sel_I[3].z ;
 wire \zbuf_bus_sel_I[4].genblk1.l ;
 wire \zbuf_bus_sel_I[4].z ;

 sky130_fd_sc_hd__clkinv_1 _18_ (.A(addr[1]),
    .Y(_00_));
 sky130_fd_sc_hd__clkinv_1 _19_ (.A(spine_iw[8]),
    .Y(_01_));
 sky130_fd_sc_hd__clkinv_1 _20_ (.A(spine_iw[9]),
    .Y(_02_));
 sky130_fd_sc_hd__clkinv_1 _21_ (.A(addr[3]),
    .Y(_03_));
 sky130_fd_sc_hd__clkinv_1 _22_ (.A(spine_iw[10]),
    .Y(_04_));
 sky130_fd_sc_hd__clkinv_1 _23_ (.A(addr[4]),
    .Y(_05_));
 sky130_fd_sc_hd__clkinv_1 _24_ (.A(\zbuf_bus_sel_I[0].z ),
    .Y(_06_));
 sky130_fd_sc_hd__clkinv_1 _25_ (.A(\zbuf_bus_sel_I[1].z ),
    .Y(_07_));
 sky130_fd_sc_hd__nor3_1 _26_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C(\zbuf_bus_sel_I[3].z ),
    .Y(\col[0].genblk1.tbuf_row_ena_I.t ));
 sky130_fd_sc_hd__nor3b_1 _27_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[3].z ),
    .C_N(\zbuf_bus_sel_I[2].z ),
    .Y(\col[2].genblk1.tbuf_row_ena_I.t ));
 sky130_fd_sc_hd__nor3b_1 _28_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C_N(\zbuf_bus_sel_I[3].z ),
    .Y(\col[4].genblk1.tbuf_row_ena_I.t ));
 sky130_fd_sc_hd__and3b_1 _29_ (.A_N(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C(\zbuf_bus_sel_I[3].z ),
    .X(\col[6].genblk1.tbuf_row_ena_I.t ));
 sky130_fd_sc_hd__xnor2_1 _30_ (.A(addr[0]),
    .B(spine_iw[6]),
    .Y(_08_));
 sky130_fd_sc_hd__o221a_1 _31_ (.A1(addr[2]),
    .A2(_02_),
    .B1(_05_),
    .B2(spine_iw[11]),
    .C1(_08_),
    .X(_09_));
 sky130_fd_sc_hd__a222oi_1 _32_ (.A1(addr[1]),
    .A2(_01_),
    .B1(_03_),
    .B2(spine_iw[10]),
    .C1(_05_),
    .C2(spine_iw[11]),
    .Y(_10_));
 sky130_fd_sc_hd__a222oi_1 _33_ (.A1(_00_),
    .A2(spine_iw[8]),
    .B1(addr[2]),
    .B2(_02_),
    .C1(addr[3]),
    .C2(_04_),
    .Y(_11_));
 sky130_fd_sc_hd__and3_1 _34_ (.A(_09_),
    .B(_10_),
    .C(_11_),
    .X(\tbuf_row_ena_I.t ));
 sky130_fd_sc_hd__nand2_1 _35_ (.A(\zbuf_bus_ena_I.z ),
    .B(\col[0].genblk1.tbuf_row_ena_I.t ),
    .Y(_12_));
 sky130_fd_sc_hd__nor3_1 _36_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_12_),
    .Y(\col[0].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _37_ (.A(_06_),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_12_),
    .Y(\col[0].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nand3_1 _38_ (.A(\zbuf_bus_ena_I.z ),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(\col[0].genblk1.tbuf_row_ena_I.t ),
    .Y(_13_));
 sky130_fd_sc_hd__nor2_1 _39_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(_13_),
    .Y(\col[1].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor2_1 _40_ (.A(_06_),
    .B(_13_),
    .Y(\col[1].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nor4bb_1 _41_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[3].z ),
    .C_N(\zbuf_bus_ena_I.z ),
    .D_N(\zbuf_bus_sel_I[2].z ),
    .Y(_14_));
 sky130_fd_sc_hd__and3_1 _42_ (.A(_06_),
    .B(_07_),
    .C(_14_),
    .X(\col[2].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__and3_1 _43_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(_07_),
    .C(_14_),
    .X(\col[2].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nand2_1 _44_ (.A(\zbuf_bus_sel_I[1].z ),
    .B(_14_),
    .Y(_15_));
 sky130_fd_sc_hd__nor2_1 _45_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(_15_),
    .Y(\col[3].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor2_1 _46_ (.A(_06_),
    .B(_15_),
    .Y(\col[3].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nand2_1 _47_ (.A(\zbuf_bus_ena_I.z ),
    .B(\col[4].genblk1.tbuf_row_ena_I.t ),
    .Y(_16_));
 sky130_fd_sc_hd__nor3_1 _48_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_16_),
    .Y(\col[4].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _49_ (.A(_06_),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_16_),
    .Y(\col[4].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _50_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(_07_),
    .C(_16_),
    .Y(\col[5].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _51_ (.A(_06_),
    .B(_07_),
    .C(_16_),
    .Y(\col[5].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nand2_1 _52_ (.A(\zbuf_bus_ena_I.z ),
    .B(\col[6].genblk1.tbuf_row_ena_I.t ),
    .Y(_17_));
 sky130_fd_sc_hd__nor3_1 _53_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_17_),
    .Y(\col[6].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _54_ (.A(_06_),
    .B(\zbuf_bus_sel_I[1].z ),
    .C(_17_),
    .Y(\col[6].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _55_ (.A(\zbuf_bus_sel_I[0].z ),
    .B(_07_),
    .C(_17_),
    .Y(\col[7].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__nor3_1 _56_ (.A(_06_),
    .B(_07_),
    .C(_17_),
    .Y(\col[7].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[0]),
    .A1(um_ow[24]),
    .A2(um_ow[48]),
    .A3(um_ow[72]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[10]),
    .A1(um_ow[34]),
    .A2(um_ow[58]),
    .A3(um_ow[82]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[11]),
    .A1(um_ow[35]),
    .A2(um_ow[59]),
    .A3(um_ow[83]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[12]),
    .A1(um_ow[36]),
    .A2(um_ow[60]),
    .A3(um_ow[84]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[13]),
    .A1(um_ow[37]),
    .A2(um_ow[61]),
    .A3(um_ow[85]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[14]),
    .A1(um_ow[38]),
    .A2(um_ow[62]),
    .A3(um_ow[86]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[15]),
    .A1(um_ow[39]),
    .A2(um_ow[63]),
    .A3(um_ow[87]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[16]),
    .A1(um_ow[40]),
    .A2(um_ow[64]),
    .A3(um_ow[88]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[17]),
    .A1(um_ow[41]),
    .A2(um_ow[65]),
    .A3(um_ow[89]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[18]),
    .A1(um_ow[42]),
    .A2(um_ow[66]),
    .A3(um_ow[90]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[19]),
    .A1(um_ow[43]),
    .A2(um_ow[67]),
    .A3(um_ow[91]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[1]),
    .A1(um_ow[25]),
    .A2(um_ow[49]),
    .A3(um_ow[73]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[20]),
    .A1(um_ow[44]),
    .A2(um_ow[68]),
    .A3(um_ow[92]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[21]),
    .A1(um_ow[45]),
    .A2(um_ow[69]),
    .A3(um_ow[93]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[22]),
    .A1(um_ow[46]),
    .A2(um_ow[70]),
    .A3(um_ow[94]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[23]),
    .A1(um_ow[47]),
    .A2(um_ow[71]),
    .A3(um_ow[95]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[2]),
    .A1(um_ow[26]),
    .A2(um_ow[50]),
    .A3(um_ow[74]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[3]),
    .A1(um_ow[27]),
    .A2(um_ow[51]),
    .A3(um_ow[75]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[4]),
    .A1(um_ow[28]),
    .A2(um_ow[52]),
    .A3(um_ow[76]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[5]),
    .A1(um_ow[29]),
    .A2(um_ow[53]),
    .A3(um_ow[77]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[6]),
    .A1(um_ow[30]),
    .A2(um_ow[54]),
    .A3(um_ow[78]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[7]),
    .A1(um_ow[31]),
    .A2(um_ow[55]),
    .A3(um_ow[79]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[8]),
    .A1(um_ow[32]),
    .A2(um_ow[56]),
    .A3(um_ow[80]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[0].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[9]),
    .A1(um_ow[33]),
    .A2(um_ow[57]),
    .A3(um_ow[81]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[0].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__inv_4 \col[0].genblk1.tbuf_row_ena_I.cell0_I  (.A(\col[0].genblk1.tbuf_row_ena_I.t ),
    .Y(\col[0].genblk1.tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[0].cell0_I  (.A(\col[0].genblk1.mux4_I[0].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[10].cell0_I  (.A(\col[0].genblk1.mux4_I[10].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[11].cell0_I  (.A(\col[0].genblk1.mux4_I[11].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[12].cell0_I  (.A(\col[0].genblk1.mux4_I[12].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[13].cell0_I  (.A(\col[0].genblk1.mux4_I[13].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[14].cell0_I  (.A(\col[0].genblk1.mux4_I[14].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[15].cell0_I  (.A(\col[0].genblk1.mux4_I[15].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[16].cell0_I  (.A(\col[0].genblk1.mux4_I[16].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[17].cell0_I  (.A(\col[0].genblk1.mux4_I[17].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[18].cell0_I  (.A(\col[0].genblk1.mux4_I[18].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[19].cell0_I  (.A(\col[0].genblk1.mux4_I[19].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[1].cell0_I  (.A(\col[0].genblk1.mux4_I[1].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[20].cell0_I  (.A(\col[0].genblk1.mux4_I[20].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[21].cell0_I  (.A(\col[0].genblk1.mux4_I[21].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[22].cell0_I  (.A(\col[0].genblk1.mux4_I[22].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[23].cell0_I  (.A(\col[0].genblk1.mux4_I[23].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[2].cell0_I  (.A(\col[0].genblk1.mux4_I[2].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[3].cell0_I  (.A(\col[0].genblk1.mux4_I[3].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[4].cell0_I  (.A(\col[0].genblk1.mux4_I[4].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[5].cell0_I  (.A(\col[0].genblk1.mux4_I[5].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[6].cell0_I  (.A(\col[0].genblk1.mux4_I[6].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[7].cell0_I  (.A(\col[0].genblk1.mux4_I[7].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[8].cell0_I  (.A(\col[0].genblk1.mux4_I[8].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \col[0].genblk1.tbuf_spine_ow_I[9].cell0_I  (.A(\col[0].genblk1.mux4_I[9].x ),
    .TE_B(\col[0].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[0].tie_bot_I.cell_I  (.HI(\col[0].tie_bot_I.hi ),
    .LO(\col[0].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[0].tie_top_I.cell_I  (.HI(\col[0].tie_top_I.hi ),
    .LO(\col[0].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[0].zbuf_bot_ena_I.e ),
    .X(\col[0].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[0].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[0].zbuf_top_ena_I.e ),
    .X(\col[0].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[1].tie_bot_I.cell_I  (.HI(\col[1].tie_bot_I.hi ),
    .LO(\col[1].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[1].tie_top_I.cell_I  (.HI(\col[1].tie_top_I.hi ),
    .LO(\col[1].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[1].zbuf_bot_ena_I.e ),
    .X(\col[1].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[1].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[1].zbuf_top_ena_I.e ),
    .X(\col[1].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[96]),
    .A1(um_ow[120]),
    .A2(um_ow[144]),
    .A3(um_ow[168]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[106]),
    .A1(um_ow[130]),
    .A2(um_ow[154]),
    .A3(um_ow[178]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[107]),
    .A1(um_ow[131]),
    .A2(um_ow[155]),
    .A3(um_ow[179]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[108]),
    .A1(um_ow[132]),
    .A2(um_ow[156]),
    .A3(um_ow[180]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[109]),
    .A1(um_ow[133]),
    .A2(um_ow[157]),
    .A3(um_ow[181]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[110]),
    .A1(um_ow[134]),
    .A2(um_ow[158]),
    .A3(um_ow[182]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[111]),
    .A1(um_ow[135]),
    .A2(um_ow[159]),
    .A3(um_ow[183]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[112]),
    .A1(um_ow[136]),
    .A2(um_ow[160]),
    .A3(um_ow[184]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[113]),
    .A1(um_ow[137]),
    .A2(um_ow[161]),
    .A3(um_ow[185]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[114]),
    .A1(um_ow[138]),
    .A2(um_ow[162]),
    .A3(um_ow[186]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[115]),
    .A1(um_ow[139]),
    .A2(um_ow[163]),
    .A3(um_ow[187]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[97]),
    .A1(um_ow[121]),
    .A2(um_ow[145]),
    .A3(um_ow[169]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[116]),
    .A1(um_ow[140]),
    .A2(um_ow[164]),
    .A3(um_ow[188]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[117]),
    .A1(um_ow[141]),
    .A2(um_ow[165]),
    .A3(um_ow[189]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[118]),
    .A1(um_ow[142]),
    .A2(um_ow[166]),
    .A3(um_ow[190]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[119]),
    .A1(um_ow[143]),
    .A2(um_ow[167]),
    .A3(um_ow[191]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[98]),
    .A1(um_ow[122]),
    .A2(um_ow[146]),
    .A3(um_ow[170]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[99]),
    .A1(um_ow[123]),
    .A2(um_ow[147]),
    .A3(um_ow[171]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[100]),
    .A1(um_ow[124]),
    .A2(um_ow[148]),
    .A3(um_ow[172]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[101]),
    .A1(um_ow[125]),
    .A2(um_ow[149]),
    .A3(um_ow[173]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[102]),
    .A1(um_ow[126]),
    .A2(um_ow[150]),
    .A3(um_ow[174]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[103]),
    .A1(um_ow[127]),
    .A2(um_ow[151]),
    .A3(um_ow[175]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[104]),
    .A1(um_ow[128]),
    .A2(um_ow[152]),
    .A3(um_ow[176]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[105]),
    .A1(um_ow[129]),
    .A2(um_ow[153]),
    .A3(um_ow[177]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[2].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__inv_4 \col[2].genblk1.tbuf_row_ena_I.cell0_I  (.A(\col[2].genblk1.tbuf_row_ena_I.t ),
    .Y(\col[2].genblk1.tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[0].cell0_I  (.A(\col[2].genblk1.mux4_I[0].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[10].cell0_I  (.A(\col[2].genblk1.mux4_I[10].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[11].cell0_I  (.A(\col[2].genblk1.mux4_I[11].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[12].cell0_I  (.A(\col[2].genblk1.mux4_I[12].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[13].cell0_I  (.A(\col[2].genblk1.mux4_I[13].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[14].cell0_I  (.A(\col[2].genblk1.mux4_I[14].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[15].cell0_I  (.A(\col[2].genblk1.mux4_I[15].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[16].cell0_I  (.A(\col[2].genblk1.mux4_I[16].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[17].cell0_I  (.A(\col[2].genblk1.mux4_I[17].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[18].cell0_I  (.A(\col[2].genblk1.mux4_I[18].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[19].cell0_I  (.A(\col[2].genblk1.mux4_I[19].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[1].cell0_I  (.A(\col[2].genblk1.mux4_I[1].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[20].cell0_I  (.A(\col[2].genblk1.mux4_I[20].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[21].cell0_I  (.A(\col[2].genblk1.mux4_I[21].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[22].cell0_I  (.A(\col[2].genblk1.mux4_I[22].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[23].cell0_I  (.A(\col[2].genblk1.mux4_I[23].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[2].cell0_I  (.A(\col[2].genblk1.mux4_I[2].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[3].cell0_I  (.A(\col[2].genblk1.mux4_I[3].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[4].cell0_I  (.A(\col[2].genblk1.mux4_I[4].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[5].cell0_I  (.A(\col[2].genblk1.mux4_I[5].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[6].cell0_I  (.A(\col[2].genblk1.mux4_I[6].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[7].cell0_I  (.A(\col[2].genblk1.mux4_I[7].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[8].cell0_I  (.A(\col[2].genblk1.mux4_I[8].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \col[2].genblk1.tbuf_spine_ow_I[9].cell0_I  (.A(\col[2].genblk1.mux4_I[9].x ),
    .TE_B(\col[2].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[2].tie_bot_I.cell_I  (.HI(\col[2].tie_bot_I.hi ),
    .LO(\col[2].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[2].tie_top_I.cell_I  (.HI(\col[2].tie_top_I.hi ),
    .LO(\col[2].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[2].zbuf_bot_ena_I.e ),
    .X(\col[2].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[2].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[2].zbuf_top_ena_I.e ),
    .X(\col[2].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[3].tie_bot_I.cell_I  (.HI(\col[3].tie_bot_I.hi ),
    .LO(\col[3].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[3].tie_top_I.cell_I  (.HI(\col[3].tie_top_I.hi ),
    .LO(\col[3].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[3].zbuf_bot_ena_I.e ),
    .X(\col[3].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[3].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[3].zbuf_top_ena_I.e ),
    .X(\col[3].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[192]),
    .A1(um_ow[216]),
    .A2(um_ow[240]),
    .A3(um_ow[264]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[202]),
    .A1(um_ow[226]),
    .A2(um_ow[250]),
    .A3(um_ow[274]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[203]),
    .A1(um_ow[227]),
    .A2(um_ow[251]),
    .A3(um_ow[275]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[204]),
    .A1(um_ow[228]),
    .A2(um_ow[252]),
    .A3(um_ow[276]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[205]),
    .A1(um_ow[229]),
    .A2(um_ow[253]),
    .A3(um_ow[277]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[206]),
    .A1(um_ow[230]),
    .A2(um_ow[254]),
    .A3(um_ow[278]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[207]),
    .A1(um_ow[231]),
    .A2(um_ow[255]),
    .A3(um_ow[279]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[208]),
    .A1(um_ow[232]),
    .A2(um_ow[256]),
    .A3(um_ow[280]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[209]),
    .A1(um_ow[233]),
    .A2(um_ow[257]),
    .A3(um_ow[281]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[210]),
    .A1(um_ow[234]),
    .A2(um_ow[258]),
    .A3(um_ow[282]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[211]),
    .A1(um_ow[235]),
    .A2(um_ow[259]),
    .A3(um_ow[283]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[193]),
    .A1(um_ow[217]),
    .A2(um_ow[241]),
    .A3(um_ow[265]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[212]),
    .A1(um_ow[236]),
    .A2(um_ow[260]),
    .A3(um_ow[284]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[213]),
    .A1(um_ow[237]),
    .A2(um_ow[261]),
    .A3(um_ow[285]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[214]),
    .A1(um_ow[238]),
    .A2(um_ow[262]),
    .A3(um_ow[286]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[215]),
    .A1(um_ow[239]),
    .A2(um_ow[263]),
    .A3(um_ow[287]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[194]),
    .A1(um_ow[218]),
    .A2(um_ow[242]),
    .A3(um_ow[266]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[195]),
    .A1(um_ow[219]),
    .A2(um_ow[243]),
    .A3(um_ow[267]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[196]),
    .A1(um_ow[220]),
    .A2(um_ow[244]),
    .A3(um_ow[268]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[197]),
    .A1(um_ow[221]),
    .A2(um_ow[245]),
    .A3(um_ow[269]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[198]),
    .A1(um_ow[222]),
    .A2(um_ow[246]),
    .A3(um_ow[270]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[199]),
    .A1(um_ow[223]),
    .A2(um_ow[247]),
    .A3(um_ow[271]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[200]),
    .A1(um_ow[224]),
    .A2(um_ow[248]),
    .A3(um_ow[272]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[201]),
    .A1(um_ow[225]),
    .A2(um_ow[249]),
    .A3(um_ow[273]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[4].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__inv_4 \col[4].genblk1.tbuf_row_ena_I.cell0_I  (.A(\col[4].genblk1.tbuf_row_ena_I.t ),
    .Y(\col[4].genblk1.tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[0].cell0_I  (.A(\col[4].genblk1.mux4_I[0].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[10].cell0_I  (.A(\col[4].genblk1.mux4_I[10].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[11].cell0_I  (.A(\col[4].genblk1.mux4_I[11].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[12].cell0_I  (.A(\col[4].genblk1.mux4_I[12].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[13].cell0_I  (.A(\col[4].genblk1.mux4_I[13].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[14].cell0_I  (.A(\col[4].genblk1.mux4_I[14].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[15].cell0_I  (.A(\col[4].genblk1.mux4_I[15].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[16].cell0_I  (.A(\col[4].genblk1.mux4_I[16].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[17].cell0_I  (.A(\col[4].genblk1.mux4_I[17].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[18].cell0_I  (.A(\col[4].genblk1.mux4_I[18].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[19].cell0_I  (.A(\col[4].genblk1.mux4_I[19].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[1].cell0_I  (.A(\col[4].genblk1.mux4_I[1].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[20].cell0_I  (.A(\col[4].genblk1.mux4_I[20].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[21].cell0_I  (.A(\col[4].genblk1.mux4_I[21].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[22].cell0_I  (.A(\col[4].genblk1.mux4_I[22].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[23].cell0_I  (.A(\col[4].genblk1.mux4_I[23].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[2].cell0_I  (.A(\col[4].genblk1.mux4_I[2].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[3].cell0_I  (.A(\col[4].genblk1.mux4_I[3].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[4].cell0_I  (.A(\col[4].genblk1.mux4_I[4].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[5].cell0_I  (.A(\col[4].genblk1.mux4_I[5].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[6].cell0_I  (.A(\col[4].genblk1.mux4_I[6].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[7].cell0_I  (.A(\col[4].genblk1.mux4_I[7].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[8].cell0_I  (.A(\col[4].genblk1.mux4_I[8].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \col[4].genblk1.tbuf_spine_ow_I[9].cell0_I  (.A(\col[4].genblk1.mux4_I[9].x ),
    .TE_B(\col[4].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[4].tie_bot_I.cell_I  (.HI(\col[4].tie_bot_I.hi ),
    .LO(\col[4].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[4].tie_top_I.cell_I  (.HI(\col[4].tie_top_I.hi ),
    .LO(\col[4].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[4].zbuf_bot_ena_I.e ),
    .X(\col[4].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[4].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[4].zbuf_top_ena_I.e ),
    .X(\col[4].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[5].tie_bot_I.cell_I  (.HI(\col[5].tie_bot_I.hi ),
    .LO(\col[5].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[5].tie_top_I.cell_I  (.HI(\col[5].tie_top_I.hi ),
    .LO(\col[5].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[5].zbuf_bot_ena_I.e ),
    .X(\col[5].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[5].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[5].zbuf_top_ena_I.e ),
    .X(\col[5].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[288]),
    .A1(um_ow[312]),
    .A2(um_ow[336]),
    .A3(um_ow[360]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[298]),
    .A1(um_ow[322]),
    .A2(um_ow[346]),
    .A3(um_ow[370]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[299]),
    .A1(um_ow[323]),
    .A2(um_ow[347]),
    .A3(um_ow[371]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[300]),
    .A1(um_ow[324]),
    .A2(um_ow[348]),
    .A3(um_ow[372]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[301]),
    .A1(um_ow[325]),
    .A2(um_ow[349]),
    .A3(um_ow[373]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[302]),
    .A1(um_ow[326]),
    .A2(um_ow[350]),
    .A3(um_ow[374]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[303]),
    .A1(um_ow[327]),
    .A2(um_ow[351]),
    .A3(um_ow[375]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[304]),
    .A1(um_ow[328]),
    .A2(um_ow[352]),
    .A3(um_ow[376]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[305]),
    .A1(um_ow[329]),
    .A2(um_ow[353]),
    .A3(um_ow[377]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[306]),
    .A1(um_ow[330]),
    .A2(um_ow[354]),
    .A3(um_ow[378]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[307]),
    .A1(um_ow[331]),
    .A2(um_ow[355]),
    .A3(um_ow[379]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[289]),
    .A1(um_ow[313]),
    .A2(um_ow[337]),
    .A3(um_ow[361]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[308]),
    .A1(um_ow[332]),
    .A2(um_ow[356]),
    .A3(um_ow[380]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[309]),
    .A1(um_ow[333]),
    .A2(um_ow[357]),
    .A3(um_ow[381]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[310]),
    .A1(um_ow[334]),
    .A2(um_ow[358]),
    .A3(um_ow[382]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[311]),
    .A1(um_ow[335]),
    .A2(um_ow[359]),
    .A3(um_ow[383]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[290]),
    .A1(um_ow[314]),
    .A2(um_ow[338]),
    .A3(um_ow[362]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[291]),
    .A1(um_ow[315]),
    .A2(um_ow[339]),
    .A3(um_ow[363]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[292]),
    .A1(um_ow[316]),
    .A2(um_ow[340]),
    .A3(um_ow[364]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[293]),
    .A1(um_ow[317]),
    .A2(um_ow[341]),
    .A3(um_ow[365]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[294]),
    .A1(um_ow[318]),
    .A2(um_ow[342]),
    .A3(um_ow[366]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[295]),
    .A1(um_ow[319]),
    .A2(um_ow[343]),
    .A3(um_ow[367]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[296]),
    .A1(um_ow[320]),
    .A2(um_ow[344]),
    .A3(um_ow[368]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[297]),
    .A1(um_ow[321]),
    .A2(um_ow[345]),
    .A3(um_ow[369]),
    .S0(\zbuf_bus_sel_I[0].z ),
    .S1(\zbuf_bus_sel_I[1].z ),
    .X(\col[6].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__inv_4 \col[6].genblk1.tbuf_row_ena_I.cell0_I  (.A(\col[6].genblk1.tbuf_row_ena_I.t ),
    .Y(\col[6].genblk1.tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[0].cell0_I  (.A(\col[6].genblk1.mux4_I[0].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[10].cell0_I  (.A(\col[6].genblk1.mux4_I[10].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[11].cell0_I  (.A(\col[6].genblk1.mux4_I[11].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[12].cell0_I  (.A(\col[6].genblk1.mux4_I[12].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[13].cell0_I  (.A(\col[6].genblk1.mux4_I[13].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[14].cell0_I  (.A(\col[6].genblk1.mux4_I[14].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[15].cell0_I  (.A(\col[6].genblk1.mux4_I[15].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[16].cell0_I  (.A(\col[6].genblk1.mux4_I[16].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[17].cell0_I  (.A(\col[6].genblk1.mux4_I[17].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[18].cell0_I  (.A(\col[6].genblk1.mux4_I[18].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[19].cell0_I  (.A(\col[6].genblk1.mux4_I[19].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[1].cell0_I  (.A(\col[6].genblk1.mux4_I[1].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[20].cell0_I  (.A(\col[6].genblk1.mux4_I[20].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[21].cell0_I  (.A(\col[6].genblk1.mux4_I[21].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[22].cell0_I  (.A(\col[6].genblk1.mux4_I[22].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[23].cell0_I  (.A(\col[6].genblk1.mux4_I[23].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[2].cell0_I  (.A(\col[6].genblk1.mux4_I[2].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[3].cell0_I  (.A(\col[6].genblk1.mux4_I[3].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[4].cell0_I  (.A(\col[6].genblk1.mux4_I[4].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[5].cell0_I  (.A(\col[6].genblk1.mux4_I[5].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[6].cell0_I  (.A(\col[6].genblk1.mux4_I[6].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[7].cell0_I  (.A(\col[6].genblk1.mux4_I[7].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[8].cell0_I  (.A(\col[6].genblk1.mux4_I[8].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \col[6].genblk1.tbuf_spine_ow_I[9].cell0_I  (.A(\col[6].genblk1.mux4_I[9].x ),
    .TE_B(\col[6].genblk1.tbuf_row_ena_I.tx ),
    .Z(\col[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[6].tie_bot_I.cell_I  (.HI(\col[6].tie_bot_I.hi ),
    .LO(\col[6].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[6].tie_top_I.cell_I  (.HI(\col[6].tie_top_I.hi ),
    .LO(\col[6].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[6].zbuf_bot_ena_I.e ),
    .X(\col[6].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[6].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[6].zbuf_top_ena_I.e ),
    .X(\col[6].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__conb_1 \col[7].tie_bot_I.cell_I  (.HI(\col[7].tie_bot_I.hi ),
    .LO(\col[7].tie_bot_I.lo ));
 sky130_fd_sc_hd__conb_1 \col[7].tie_top_I.cell_I  (.HI(\col[7].tie_top_I.hi ),
    .LO(\col[7].tie_top_I.lo ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[7].zbuf_bot_ena_I.e ),
    .X(\col[7].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \col[7].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .B(\col[7].zbuf_top_ena_I.e ),
    .X(\col[7].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__inv_4 \tbuf_row_ena_I.cell0_I  (.A(\tbuf_row_ena_I.t ),
    .Y(\tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[0].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[0].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[10].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[10].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[11].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[11].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[12].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[12].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[13].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[13].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[14].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[14].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[15].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[15].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[16].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[16].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[17].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[17].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[18].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[18].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[19].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[19].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[1].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[1].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[20].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[20].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[21].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[21].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[22].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[22].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[23].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[23].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[2].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[2].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[3].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[3].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[4].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[4].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[5].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[5].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[6].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[6].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[7].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[7].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[8].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[8].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[9].cell0_I  (.A(\col[0].genblk1.tbuf_spine_ow_I[9].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \tie_I.cell_I  (.HI(k_one),
    .LO(k_zero));
 sky130_fd_sc_hd__conb_1 \tie_spine_guard_I[0].cell_I  (.HI(\tie_spine_guard_I[0].hi ),
    .LO(\tie_spine_guard_I[0].lo ));
 sky130_fd_sc_hd__conb_1 \tie_spine_guard_I[1].cell_I  (.HI(\tie_spine_guard_I[1].hi ),
    .LO(\tie_spine_guard_I[1].lo ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_ena_I.genblk1.cell0_I  (.A(spine_iw[1]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_ena_I.genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_ena_I.genblk1.cell1_I  (.A(\zbuf_bus_ena_I.genblk1.l ),
    .X(\zbuf_bus_ena_I.z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[0].genblk1.cell0_I  (.A(spine_iw[12]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[0].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[0].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[10].genblk1.cell0_I  (.A(spine_iw[22]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[10].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[10].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[10].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[11].genblk1.cell0_I  (.A(spine_iw[23]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[11].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[11].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[11].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[12].genblk1.cell0_I  (.A(spine_iw[24]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[12].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[12].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[12].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[13].genblk1.cell0_I  (.A(spine_iw[25]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[13].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[13].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[13].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[14].genblk1.cell0_I  (.A(spine_iw[26]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[14].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[14].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[14].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[15].genblk1.cell0_I  (.A(spine_iw[27]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[15].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[15].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[15].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[16].genblk1.cell0_I  (.A(spine_iw[28]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[16].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[16].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[16].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[17].genblk1.cell0_I  (.A(spine_iw[29]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[17].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[17].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[17].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[1].genblk1.cell0_I  (.A(spine_iw[13]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[1].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[1].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[2].genblk1.cell0_I  (.A(spine_iw[14]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[2].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[2].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[3].genblk1.cell0_I  (.A(spine_iw[15]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[3].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[3].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[4].genblk1.cell0_I  (.A(spine_iw[16]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[4].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[4].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[5].genblk1.cell0_I  (.A(spine_iw[17]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[5].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[5].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[6].genblk1.cell0_I  (.A(spine_iw[18]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[6].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[6].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[7].genblk1.cell0_I  (.A(spine_iw[19]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[7].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[7].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[8].genblk1.cell0_I  (.A(spine_iw[20]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[8].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[8].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[9].genblk1.cell0_I  (.A(spine_iw[21]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_iw_I[9].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[9].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[9].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[0].genblk1.cell0_I  (.A(spine_iw[7]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_sel_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[0].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[0].genblk1.l ),
    .X(\zbuf_bus_sel_I[0].z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[1].genblk1.cell0_I  (.A(spine_iw[2]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_sel_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[1].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[1].genblk1.l ),
    .X(\zbuf_bus_sel_I[1].z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[2].genblk1.cell0_I  (.A(spine_iw[3]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_sel_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[2].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[2].genblk1.l ),
    .X(\zbuf_bus_sel_I[2].z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[3].genblk1.cell0_I  (.A(spine_iw[4]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_sel_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[3].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[3].genblk1.l ),
    .X(\zbuf_bus_sel_I[3].z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[4].genblk1.cell0_I  (.A(spine_iw[5]),
    .B(\tbuf_row_ena_I.t ),
    .X(\zbuf_bus_sel_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[4].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[4].genblk1.l ),
    .X(\zbuf_bus_sel_I[4].z ));
 sky130_fd_sc_hd__conb_1 TIE_ONE_one_ (.HI(one_));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\col[1].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\col[2].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\col[6].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(\col[6].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(\col[6].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(spine_iw[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(spine_iw[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(spine_iw[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(um_ow[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(um_ow[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(um_ow[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(um_ow[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(um_ow[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(um_ow[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(um_ow[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(um_ow[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(um_ow[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(um_ow[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(um_ow[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(um_ow[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(um_ow[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(um_ow[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(um_ow[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(um_ow[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(um_ow[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(um_ow[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(um_ow[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(um_ow[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(um_ow[124]));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(um_ow[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(um_ow[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(um_ow[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(um_ow[128]));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(um_ow[129]));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(um_ow[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(um_ow[131]));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(um_ow[132]));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(um_ow[133]));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(um_ow[135]));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(um_ow[137]));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(um_ow[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(um_ow[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(um_ow[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(um_ow[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(um_ow[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(um_ow[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(um_ow[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(um_ow[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(um_ow[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(um_ow[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(um_ow[240]));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(um_ow[241]));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(um_ow[242]));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(um_ow[243]));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(um_ow[244]));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(um_ow[245]));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(um_ow[246]));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(um_ow[247]));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(um_ow[248]));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(um_ow[249]));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(um_ow[250]));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(um_ow[251]));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(um_ow[252]));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(um_ow[253]));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(um_ow[254]));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(um_ow[255]));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(um_ow[257]));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(um_ow[258]));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(um_ow[259]));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(um_ow[260]));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(um_ow[261]));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(um_ow[263]));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(um_ow[269]));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(um_ow[270]));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(um_ow[271]));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(um_ow[272]));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(um_ow[273]));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(um_ow[274]));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(um_ow[275]));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(um_ow[278]));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(um_ow[279]));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(um_ow[281]));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(um_ow[283]));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(um_ow[284]));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(um_ow[285]));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(um_ow[286]));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(um_ow[287]));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(um_ow[336]));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(um_ow[337]));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(um_ow[338]));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(um_ow[339]));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(um_ow[340]));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(um_ow[341]));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(um_ow[342]));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(um_ow[343]));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(um_ow[344]));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(um_ow[345]));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(um_ow[346]));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(um_ow[347]));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(um_ow[348]));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(um_ow[349]));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(um_ow[350]));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(um_ow[351]));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(um_ow[352]));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(um_ow[353]));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(um_ow[354]));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(um_ow[355]));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(um_ow[356]));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(um_ow[357]));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(um_ow[358]));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(um_ow[359]));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(um_ow[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(um_ow[360]));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(um_ow[370]));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(um_ow[371]));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(um_ow[373]));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(um_ow[376]));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(um_ow[380]));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(um_ow[381]));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(um_ow[382]));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(um_ow[383]));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(um_ow[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(um_ow[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(um_ow[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(um_ow[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(um_ow[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(um_ow[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(um_ow[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(um_ow[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(um_ow[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(um_ow[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(um_ow[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(um_ow[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(um_ow[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(um_ow[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(um_ow[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(um_ow[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(um_ow[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\col[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\col[0].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(um_ow[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(um_ow[136]));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(um_ow[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(um_ow[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(um_ow[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(um_ow[140]));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(um_ow[29]));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1295 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1387 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1448 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1555 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1563 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1611 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1615 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1619 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1646 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1671 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1693 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1701 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1717 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1773 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1871 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1883 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1895 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2061 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2067 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2070 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2073 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2078 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2086 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2094 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2102 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2118 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2126 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2135 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2150 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2157 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2191 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2218 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2230 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2262 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2287 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2309 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2313 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2365 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2395 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2430 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2455 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2459 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2477 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2512 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2554 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2566 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2574 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2589 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2745 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2780 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2793 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2801 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2809 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2817 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2835 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2844 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2852 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2875 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2882 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2890 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2899 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2911 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2934 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1639 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1730 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1755 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2225 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2233 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2237 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2264 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2281 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2285 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2367 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2402 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2427 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2437 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2459 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2638 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2650 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2658 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2785 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2811 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2823 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2841 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2847 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1555 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1622 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1625 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1654 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2247 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2251 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2297 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2313 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2353 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2363 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2386 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2406 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2432 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2498 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2510 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2518 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2554 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2566 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2574 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2778 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2790 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2798 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2825 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2850 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2881 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2934 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1290 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1562 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1609 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1633 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1637 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1645 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1667 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1713 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2269 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2321 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2325 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2353 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2356 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2661 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2692 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2704 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2794 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2806 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2818 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2826 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2850 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2862 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2921 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2927 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1646 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1655 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1876 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2330 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2342 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2350 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2406 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2421 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2429 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2433 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2460 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2498 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2510 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2518 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2554 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2566 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2574 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2645 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2676 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2772 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2881 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2934 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1585 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1639 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1678 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1682 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2281 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2319 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2325 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2333 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2356 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2360 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2418 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2897 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2909 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2925 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1544 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1573 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1585 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1588 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1619 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1646 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1654 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2295 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2297 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2321 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2374 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2378 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2403 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2550 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2562 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2574 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2930 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1527 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1590 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1601 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1650 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1656 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1675 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1687 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2841 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2845 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2858 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2866 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2897 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1628 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1636 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1640 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1663 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2208 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2216 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2228 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2813 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2848 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2857 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2909 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2934 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1633 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2437 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2449 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2457 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2530 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2841 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2853 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2895 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2929 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1649 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1655 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1664 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2489 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2869 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2905 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2935 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2461 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2473 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2493 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2507 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2514 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2520 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2897 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2909 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2915 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2933 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1605 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1631 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1635 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1671 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2911 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2934 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1634 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1646 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2897 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2909 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1420 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1428 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1436 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1713 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1797 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1803 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2071 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2073 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2079 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2086 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2094 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2100 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2107 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2119 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2153 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2160 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2168 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2176 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2433 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2507 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2519 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2521 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2531 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2539 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2547 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2563 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2813 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2827 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2835 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2842 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2854 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2881 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2901 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2909 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2913 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2935 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1458 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1462 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1671 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1675 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1683 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1692 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1701 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1715 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1719 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1725 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1729 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1741 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1757 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1816 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1821 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1825 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1857 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1865 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1871 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2025 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2033 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2038 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2045 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2053 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2062 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2078 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2082 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2086 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2094 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2098 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2119 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2126 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2142 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2150 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2154 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2191 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2199 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2225 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2393 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2405 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2416 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2424 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2432 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2449 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2453 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2457 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2465 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2469 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2481 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2489 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2505 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2513 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2521 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2529 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2537 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2545 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2561 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2565 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2771 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2779 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2782 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2786 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2794 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2802 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2818 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2822 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2826 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2834 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2838 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2842 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2850 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2867 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2875 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2891 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2899 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2907 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2926 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2930 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2917 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2925 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2932 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2936 ();
 assign um_k_zero[0] = \col[0].tie_bot_I.lo ;
 assign um_k_zero[1] = \col[0].tie_top_I.lo ;
 assign um_ena[0] = \col[0].zbuf_bot_ena_I.z ;
 assign um_iw[0] = \col[0].zbuf_bot_iw_I[0].z ;
 assign um_iw[10] = \col[0].zbuf_bot_iw_I[10].z ;
 assign um_iw[11] = \col[0].zbuf_bot_iw_I[11].z ;
 assign um_iw[12] = \col[0].zbuf_bot_iw_I[12].z ;
 assign um_iw[13] = \col[0].zbuf_bot_iw_I[13].z ;
 assign um_iw[14] = \col[0].zbuf_bot_iw_I[14].z ;
 assign um_iw[15] = \col[0].zbuf_bot_iw_I[15].z ;
 assign um_iw[16] = \col[0].zbuf_bot_iw_I[16].z ;
 assign um_iw[17] = \col[0].zbuf_bot_iw_I[17].z ;
 assign um_iw[1] = \col[0].zbuf_bot_iw_I[1].z ;
 assign um_iw[2] = \col[0].zbuf_bot_iw_I[2].z ;
 assign um_iw[3] = \col[0].zbuf_bot_iw_I[3].z ;
 assign um_iw[4] = \col[0].zbuf_bot_iw_I[4].z ;
 assign um_iw[5] = \col[0].zbuf_bot_iw_I[5].z ;
 assign um_iw[6] = \col[0].zbuf_bot_iw_I[6].z ;
 assign um_iw[7] = \col[0].zbuf_bot_iw_I[7].z ;
 assign um_iw[8] = \col[0].zbuf_bot_iw_I[8].z ;
 assign um_iw[9] = \col[0].zbuf_bot_iw_I[9].z ;
 assign um_ena[1] = \col[0].zbuf_top_ena_I.z ;
 assign um_iw[18] = \col[0].zbuf_top_iw_I[0].z ;
 assign um_iw[28] = \col[0].zbuf_top_iw_I[10].z ;
 assign um_iw[29] = \col[0].zbuf_top_iw_I[11].z ;
 assign um_iw[30] = \col[0].zbuf_top_iw_I[12].z ;
 assign um_iw[31] = \col[0].zbuf_top_iw_I[13].z ;
 assign um_iw[32] = \col[0].zbuf_top_iw_I[14].z ;
 assign um_iw[33] = \col[0].zbuf_top_iw_I[15].z ;
 assign um_iw[34] = \col[0].zbuf_top_iw_I[16].z ;
 assign um_iw[35] = \col[0].zbuf_top_iw_I[17].z ;
 assign um_iw[19] = \col[0].zbuf_top_iw_I[1].z ;
 assign um_iw[20] = \col[0].zbuf_top_iw_I[2].z ;
 assign um_iw[21] = \col[0].zbuf_top_iw_I[3].z ;
 assign um_iw[22] = \col[0].zbuf_top_iw_I[4].z ;
 assign um_iw[23] = \col[0].zbuf_top_iw_I[5].z ;
 assign um_iw[24] = \col[0].zbuf_top_iw_I[6].z ;
 assign um_iw[25] = \col[0].zbuf_top_iw_I[7].z ;
 assign um_iw[26] = \col[0].zbuf_top_iw_I[8].z ;
 assign um_iw[27] = \col[0].zbuf_top_iw_I[9].z ;
 assign um_k_zero[2] = \col[1].tie_bot_I.lo ;
 assign um_k_zero[3] = \col[1].tie_top_I.lo ;
 assign um_ena[2] = \col[1].zbuf_bot_ena_I.z ;
 assign um_iw[36] = \col[1].zbuf_bot_iw_I[0].z ;
 assign um_iw[46] = \col[1].zbuf_bot_iw_I[10].z ;
 assign um_iw[47] = \col[1].zbuf_bot_iw_I[11].z ;
 assign um_iw[48] = \col[1].zbuf_bot_iw_I[12].z ;
 assign um_iw[49] = \col[1].zbuf_bot_iw_I[13].z ;
 assign um_iw[50] = \col[1].zbuf_bot_iw_I[14].z ;
 assign um_iw[51] = \col[1].zbuf_bot_iw_I[15].z ;
 assign um_iw[52] = \col[1].zbuf_bot_iw_I[16].z ;
 assign um_iw[53] = \col[1].zbuf_bot_iw_I[17].z ;
 assign um_iw[37] = \col[1].zbuf_bot_iw_I[1].z ;
 assign um_iw[38] = \col[1].zbuf_bot_iw_I[2].z ;
 assign um_iw[39] = \col[1].zbuf_bot_iw_I[3].z ;
 assign um_iw[40] = \col[1].zbuf_bot_iw_I[4].z ;
 assign um_iw[41] = \col[1].zbuf_bot_iw_I[5].z ;
 assign um_iw[42] = \col[1].zbuf_bot_iw_I[6].z ;
 assign um_iw[43] = \col[1].zbuf_bot_iw_I[7].z ;
 assign um_iw[44] = \col[1].zbuf_bot_iw_I[8].z ;
 assign um_iw[45] = \col[1].zbuf_bot_iw_I[9].z ;
 assign um_ena[3] = \col[1].zbuf_top_ena_I.z ;
 assign um_iw[54] = \col[1].zbuf_top_iw_I[0].z ;
 assign um_iw[64] = \col[1].zbuf_top_iw_I[10].z ;
 assign um_iw[65] = \col[1].zbuf_top_iw_I[11].z ;
 assign um_iw[66] = \col[1].zbuf_top_iw_I[12].z ;
 assign um_iw[67] = \col[1].zbuf_top_iw_I[13].z ;
 assign um_iw[68] = \col[1].zbuf_top_iw_I[14].z ;
 assign um_iw[69] = \col[1].zbuf_top_iw_I[15].z ;
 assign um_iw[70] = \col[1].zbuf_top_iw_I[16].z ;
 assign um_iw[71] = \col[1].zbuf_top_iw_I[17].z ;
 assign um_iw[55] = \col[1].zbuf_top_iw_I[1].z ;
 assign um_iw[56] = \col[1].zbuf_top_iw_I[2].z ;
 assign um_iw[57] = \col[1].zbuf_top_iw_I[3].z ;
 assign um_iw[58] = \col[1].zbuf_top_iw_I[4].z ;
 assign um_iw[59] = \col[1].zbuf_top_iw_I[5].z ;
 assign um_iw[60] = \col[1].zbuf_top_iw_I[6].z ;
 assign um_iw[61] = \col[1].zbuf_top_iw_I[7].z ;
 assign um_iw[62] = \col[1].zbuf_top_iw_I[8].z ;
 assign um_iw[63] = \col[1].zbuf_top_iw_I[9].z ;
 assign um_k_zero[4] = \col[2].tie_bot_I.lo ;
 assign um_k_zero[5] = \col[2].tie_top_I.lo ;
 assign um_ena[4] = \col[2].zbuf_bot_ena_I.z ;
 assign um_iw[72] = \col[2].zbuf_bot_iw_I[0].z ;
 assign um_iw[82] = \col[2].zbuf_bot_iw_I[10].z ;
 assign um_iw[83] = \col[2].zbuf_bot_iw_I[11].z ;
 assign um_iw[84] = \col[2].zbuf_bot_iw_I[12].z ;
 assign um_iw[85] = \col[2].zbuf_bot_iw_I[13].z ;
 assign um_iw[86] = \col[2].zbuf_bot_iw_I[14].z ;
 assign um_iw[87] = \col[2].zbuf_bot_iw_I[15].z ;
 assign um_iw[88] = \col[2].zbuf_bot_iw_I[16].z ;
 assign um_iw[89] = \col[2].zbuf_bot_iw_I[17].z ;
 assign um_iw[73] = \col[2].zbuf_bot_iw_I[1].z ;
 assign um_iw[74] = \col[2].zbuf_bot_iw_I[2].z ;
 assign um_iw[75] = \col[2].zbuf_bot_iw_I[3].z ;
 assign um_iw[76] = \col[2].zbuf_bot_iw_I[4].z ;
 assign um_iw[77] = \col[2].zbuf_bot_iw_I[5].z ;
 assign um_iw[78] = \col[2].zbuf_bot_iw_I[6].z ;
 assign um_iw[79] = \col[2].zbuf_bot_iw_I[7].z ;
 assign um_iw[80] = \col[2].zbuf_bot_iw_I[8].z ;
 assign um_iw[81] = \col[2].zbuf_bot_iw_I[9].z ;
 assign um_ena[5] = \col[2].zbuf_top_ena_I.z ;
 assign um_iw[90] = \col[2].zbuf_top_iw_I[0].z ;
 assign um_iw[100] = \col[2].zbuf_top_iw_I[10].z ;
 assign um_iw[101] = \col[2].zbuf_top_iw_I[11].z ;
 assign um_iw[102] = \col[2].zbuf_top_iw_I[12].z ;
 assign um_iw[103] = \col[2].zbuf_top_iw_I[13].z ;
 assign um_iw[104] = \col[2].zbuf_top_iw_I[14].z ;
 assign um_iw[105] = \col[2].zbuf_top_iw_I[15].z ;
 assign um_iw[106] = \col[2].zbuf_top_iw_I[16].z ;
 assign um_iw[107] = \col[2].zbuf_top_iw_I[17].z ;
 assign um_iw[91] = \col[2].zbuf_top_iw_I[1].z ;
 assign um_iw[92] = \col[2].zbuf_top_iw_I[2].z ;
 assign um_iw[93] = \col[2].zbuf_top_iw_I[3].z ;
 assign um_iw[94] = \col[2].zbuf_top_iw_I[4].z ;
 assign um_iw[95] = \col[2].zbuf_top_iw_I[5].z ;
 assign um_iw[96] = \col[2].zbuf_top_iw_I[6].z ;
 assign um_iw[97] = \col[2].zbuf_top_iw_I[7].z ;
 assign um_iw[98] = \col[2].zbuf_top_iw_I[8].z ;
 assign um_iw[99] = \col[2].zbuf_top_iw_I[9].z ;
 assign um_k_zero[6] = \col[3].tie_bot_I.lo ;
 assign um_k_zero[7] = \col[3].tie_top_I.lo ;
 assign um_ena[6] = \col[3].zbuf_bot_ena_I.z ;
 assign um_iw[108] = \col[3].zbuf_bot_iw_I[0].z ;
 assign um_iw[118] = \col[3].zbuf_bot_iw_I[10].z ;
 assign um_iw[119] = \col[3].zbuf_bot_iw_I[11].z ;
 assign um_iw[120] = \col[3].zbuf_bot_iw_I[12].z ;
 assign um_iw[121] = \col[3].zbuf_bot_iw_I[13].z ;
 assign um_iw[122] = \col[3].zbuf_bot_iw_I[14].z ;
 assign um_iw[123] = \col[3].zbuf_bot_iw_I[15].z ;
 assign um_iw[124] = \col[3].zbuf_bot_iw_I[16].z ;
 assign um_iw[125] = \col[3].zbuf_bot_iw_I[17].z ;
 assign um_iw[109] = \col[3].zbuf_bot_iw_I[1].z ;
 assign um_iw[110] = \col[3].zbuf_bot_iw_I[2].z ;
 assign um_iw[111] = \col[3].zbuf_bot_iw_I[3].z ;
 assign um_iw[112] = \col[3].zbuf_bot_iw_I[4].z ;
 assign um_iw[113] = \col[3].zbuf_bot_iw_I[5].z ;
 assign um_iw[114] = \col[3].zbuf_bot_iw_I[6].z ;
 assign um_iw[115] = \col[3].zbuf_bot_iw_I[7].z ;
 assign um_iw[116] = \col[3].zbuf_bot_iw_I[8].z ;
 assign um_iw[117] = \col[3].zbuf_bot_iw_I[9].z ;
 assign um_ena[7] = \col[3].zbuf_top_ena_I.z ;
 assign um_iw[126] = \col[3].zbuf_top_iw_I[0].z ;
 assign um_iw[136] = \col[3].zbuf_top_iw_I[10].z ;
 assign um_iw[137] = \col[3].zbuf_top_iw_I[11].z ;
 assign um_iw[138] = \col[3].zbuf_top_iw_I[12].z ;
 assign um_iw[139] = \col[3].zbuf_top_iw_I[13].z ;
 assign um_iw[140] = \col[3].zbuf_top_iw_I[14].z ;
 assign um_iw[141] = \col[3].zbuf_top_iw_I[15].z ;
 assign um_iw[142] = \col[3].zbuf_top_iw_I[16].z ;
 assign um_iw[143] = \col[3].zbuf_top_iw_I[17].z ;
 assign um_iw[127] = \col[3].zbuf_top_iw_I[1].z ;
 assign um_iw[128] = \col[3].zbuf_top_iw_I[2].z ;
 assign um_iw[129] = \col[3].zbuf_top_iw_I[3].z ;
 assign um_iw[130] = \col[3].zbuf_top_iw_I[4].z ;
 assign um_iw[131] = \col[3].zbuf_top_iw_I[5].z ;
 assign um_iw[132] = \col[3].zbuf_top_iw_I[6].z ;
 assign um_iw[133] = \col[3].zbuf_top_iw_I[7].z ;
 assign um_iw[134] = \col[3].zbuf_top_iw_I[8].z ;
 assign um_iw[135] = \col[3].zbuf_top_iw_I[9].z ;
 assign um_k_zero[8] = \col[4].tie_bot_I.lo ;
 assign um_k_zero[9] = \col[4].tie_top_I.lo ;
 assign um_ena[8] = \col[4].zbuf_bot_ena_I.z ;
 assign um_iw[144] = \col[4].zbuf_bot_iw_I[0].z ;
 assign um_iw[154] = \col[4].zbuf_bot_iw_I[10].z ;
 assign um_iw[155] = \col[4].zbuf_bot_iw_I[11].z ;
 assign um_iw[156] = \col[4].zbuf_bot_iw_I[12].z ;
 assign um_iw[157] = \col[4].zbuf_bot_iw_I[13].z ;
 assign um_iw[158] = \col[4].zbuf_bot_iw_I[14].z ;
 assign um_iw[159] = \col[4].zbuf_bot_iw_I[15].z ;
 assign um_iw[160] = \col[4].zbuf_bot_iw_I[16].z ;
 assign um_iw[161] = \col[4].zbuf_bot_iw_I[17].z ;
 assign um_iw[145] = \col[4].zbuf_bot_iw_I[1].z ;
 assign um_iw[146] = \col[4].zbuf_bot_iw_I[2].z ;
 assign um_iw[147] = \col[4].zbuf_bot_iw_I[3].z ;
 assign um_iw[148] = \col[4].zbuf_bot_iw_I[4].z ;
 assign um_iw[149] = \col[4].zbuf_bot_iw_I[5].z ;
 assign um_iw[150] = \col[4].zbuf_bot_iw_I[6].z ;
 assign um_iw[151] = \col[4].zbuf_bot_iw_I[7].z ;
 assign um_iw[152] = \col[4].zbuf_bot_iw_I[8].z ;
 assign um_iw[153] = \col[4].zbuf_bot_iw_I[9].z ;
 assign um_ena[9] = \col[4].zbuf_top_ena_I.z ;
 assign um_iw[162] = \col[4].zbuf_top_iw_I[0].z ;
 assign um_iw[172] = \col[4].zbuf_top_iw_I[10].z ;
 assign um_iw[173] = \col[4].zbuf_top_iw_I[11].z ;
 assign um_iw[174] = \col[4].zbuf_top_iw_I[12].z ;
 assign um_iw[175] = \col[4].zbuf_top_iw_I[13].z ;
 assign um_iw[176] = \col[4].zbuf_top_iw_I[14].z ;
 assign um_iw[177] = \col[4].zbuf_top_iw_I[15].z ;
 assign um_iw[178] = \col[4].zbuf_top_iw_I[16].z ;
 assign um_iw[179] = \col[4].zbuf_top_iw_I[17].z ;
 assign um_iw[163] = \col[4].zbuf_top_iw_I[1].z ;
 assign um_iw[164] = \col[4].zbuf_top_iw_I[2].z ;
 assign um_iw[165] = \col[4].zbuf_top_iw_I[3].z ;
 assign um_iw[166] = \col[4].zbuf_top_iw_I[4].z ;
 assign um_iw[167] = \col[4].zbuf_top_iw_I[5].z ;
 assign um_iw[168] = \col[4].zbuf_top_iw_I[6].z ;
 assign um_iw[169] = \col[4].zbuf_top_iw_I[7].z ;
 assign um_iw[170] = \col[4].zbuf_top_iw_I[8].z ;
 assign um_iw[171] = \col[4].zbuf_top_iw_I[9].z ;
 assign um_k_zero[10] = \col[5].tie_bot_I.lo ;
 assign um_k_zero[11] = \col[5].tie_top_I.lo ;
 assign um_ena[10] = \col[5].zbuf_bot_ena_I.z ;
 assign um_iw[180] = \col[5].zbuf_bot_iw_I[0].z ;
 assign um_iw[190] = \col[5].zbuf_bot_iw_I[10].z ;
 assign um_iw[191] = \col[5].zbuf_bot_iw_I[11].z ;
 assign um_iw[192] = \col[5].zbuf_bot_iw_I[12].z ;
 assign um_iw[193] = \col[5].zbuf_bot_iw_I[13].z ;
 assign um_iw[194] = \col[5].zbuf_bot_iw_I[14].z ;
 assign um_iw[195] = \col[5].zbuf_bot_iw_I[15].z ;
 assign um_iw[196] = \col[5].zbuf_bot_iw_I[16].z ;
 assign um_iw[197] = \col[5].zbuf_bot_iw_I[17].z ;
 assign um_iw[181] = \col[5].zbuf_bot_iw_I[1].z ;
 assign um_iw[182] = \col[5].zbuf_bot_iw_I[2].z ;
 assign um_iw[183] = \col[5].zbuf_bot_iw_I[3].z ;
 assign um_iw[184] = \col[5].zbuf_bot_iw_I[4].z ;
 assign um_iw[185] = \col[5].zbuf_bot_iw_I[5].z ;
 assign um_iw[186] = \col[5].zbuf_bot_iw_I[6].z ;
 assign um_iw[187] = \col[5].zbuf_bot_iw_I[7].z ;
 assign um_iw[188] = \col[5].zbuf_bot_iw_I[8].z ;
 assign um_iw[189] = \col[5].zbuf_bot_iw_I[9].z ;
 assign um_ena[11] = \col[5].zbuf_top_ena_I.z ;
 assign um_iw[198] = \col[5].zbuf_top_iw_I[0].z ;
 assign um_iw[208] = \col[5].zbuf_top_iw_I[10].z ;
 assign um_iw[209] = \col[5].zbuf_top_iw_I[11].z ;
 assign um_iw[210] = \col[5].zbuf_top_iw_I[12].z ;
 assign um_iw[211] = \col[5].zbuf_top_iw_I[13].z ;
 assign um_iw[212] = \col[5].zbuf_top_iw_I[14].z ;
 assign um_iw[213] = \col[5].zbuf_top_iw_I[15].z ;
 assign um_iw[214] = \col[5].zbuf_top_iw_I[16].z ;
 assign um_iw[215] = \col[5].zbuf_top_iw_I[17].z ;
 assign um_iw[199] = \col[5].zbuf_top_iw_I[1].z ;
 assign um_iw[200] = \col[5].zbuf_top_iw_I[2].z ;
 assign um_iw[201] = \col[5].zbuf_top_iw_I[3].z ;
 assign um_iw[202] = \col[5].zbuf_top_iw_I[4].z ;
 assign um_iw[203] = \col[5].zbuf_top_iw_I[5].z ;
 assign um_iw[204] = \col[5].zbuf_top_iw_I[6].z ;
 assign um_iw[205] = \col[5].zbuf_top_iw_I[7].z ;
 assign um_iw[206] = \col[5].zbuf_top_iw_I[8].z ;
 assign um_iw[207] = \col[5].zbuf_top_iw_I[9].z ;
 assign um_k_zero[12] = \col[6].tie_bot_I.lo ;
 assign um_k_zero[13] = \col[6].tie_top_I.lo ;
 assign um_ena[12] = \col[6].zbuf_bot_ena_I.z ;
 assign um_iw[216] = \col[6].zbuf_bot_iw_I[0].z ;
 assign um_iw[226] = \col[6].zbuf_bot_iw_I[10].z ;
 assign um_iw[227] = \col[6].zbuf_bot_iw_I[11].z ;
 assign um_iw[228] = \col[6].zbuf_bot_iw_I[12].z ;
 assign um_iw[229] = \col[6].zbuf_bot_iw_I[13].z ;
 assign um_iw[230] = \col[6].zbuf_bot_iw_I[14].z ;
 assign um_iw[231] = \col[6].zbuf_bot_iw_I[15].z ;
 assign um_iw[232] = \col[6].zbuf_bot_iw_I[16].z ;
 assign um_iw[233] = \col[6].zbuf_bot_iw_I[17].z ;
 assign um_iw[217] = \col[6].zbuf_bot_iw_I[1].z ;
 assign um_iw[218] = \col[6].zbuf_bot_iw_I[2].z ;
 assign um_iw[219] = \col[6].zbuf_bot_iw_I[3].z ;
 assign um_iw[220] = \col[6].zbuf_bot_iw_I[4].z ;
 assign um_iw[221] = \col[6].zbuf_bot_iw_I[5].z ;
 assign um_iw[222] = \col[6].zbuf_bot_iw_I[6].z ;
 assign um_iw[223] = \col[6].zbuf_bot_iw_I[7].z ;
 assign um_iw[224] = \col[6].zbuf_bot_iw_I[8].z ;
 assign um_iw[225] = \col[6].zbuf_bot_iw_I[9].z ;
 assign um_ena[13] = \col[6].zbuf_top_ena_I.z ;
 assign um_iw[234] = \col[6].zbuf_top_iw_I[0].z ;
 assign um_iw[244] = \col[6].zbuf_top_iw_I[10].z ;
 assign um_iw[245] = \col[6].zbuf_top_iw_I[11].z ;
 assign um_iw[246] = \col[6].zbuf_top_iw_I[12].z ;
 assign um_iw[247] = \col[6].zbuf_top_iw_I[13].z ;
 assign um_iw[248] = \col[6].zbuf_top_iw_I[14].z ;
 assign um_iw[249] = \col[6].zbuf_top_iw_I[15].z ;
 assign um_iw[250] = \col[6].zbuf_top_iw_I[16].z ;
 assign um_iw[251] = \col[6].zbuf_top_iw_I[17].z ;
 assign um_iw[235] = \col[6].zbuf_top_iw_I[1].z ;
 assign um_iw[236] = \col[6].zbuf_top_iw_I[2].z ;
 assign um_iw[237] = \col[6].zbuf_top_iw_I[3].z ;
 assign um_iw[238] = \col[6].zbuf_top_iw_I[4].z ;
 assign um_iw[239] = \col[6].zbuf_top_iw_I[5].z ;
 assign um_iw[240] = \col[6].zbuf_top_iw_I[6].z ;
 assign um_iw[241] = \col[6].zbuf_top_iw_I[7].z ;
 assign um_iw[242] = \col[6].zbuf_top_iw_I[8].z ;
 assign um_iw[243] = \col[6].zbuf_top_iw_I[9].z ;
 assign um_k_zero[14] = \col[7].tie_bot_I.lo ;
 assign um_k_zero[15] = \col[7].tie_top_I.lo ;
 assign um_ena[14] = \col[7].zbuf_bot_ena_I.z ;
 assign um_iw[252] = \col[7].zbuf_bot_iw_I[0].z ;
 assign um_iw[262] = \col[7].zbuf_bot_iw_I[10].z ;
 assign um_iw[263] = \col[7].zbuf_bot_iw_I[11].z ;
 assign um_iw[264] = \col[7].zbuf_bot_iw_I[12].z ;
 assign um_iw[265] = \col[7].zbuf_bot_iw_I[13].z ;
 assign um_iw[266] = \col[7].zbuf_bot_iw_I[14].z ;
 assign um_iw[267] = \col[7].zbuf_bot_iw_I[15].z ;
 assign um_iw[268] = \col[7].zbuf_bot_iw_I[16].z ;
 assign um_iw[269] = \col[7].zbuf_bot_iw_I[17].z ;
 assign um_iw[253] = \col[7].zbuf_bot_iw_I[1].z ;
 assign um_iw[254] = \col[7].zbuf_bot_iw_I[2].z ;
 assign um_iw[255] = \col[7].zbuf_bot_iw_I[3].z ;
 assign um_iw[256] = \col[7].zbuf_bot_iw_I[4].z ;
 assign um_iw[257] = \col[7].zbuf_bot_iw_I[5].z ;
 assign um_iw[258] = \col[7].zbuf_bot_iw_I[6].z ;
 assign um_iw[259] = \col[7].zbuf_bot_iw_I[7].z ;
 assign um_iw[260] = \col[7].zbuf_bot_iw_I[8].z ;
 assign um_iw[261] = \col[7].zbuf_bot_iw_I[9].z ;
 assign um_ena[15] = \col[7].zbuf_top_ena_I.z ;
 assign um_iw[270] = \col[7].zbuf_top_iw_I[0].z ;
 assign um_iw[280] = \col[7].zbuf_top_iw_I[10].z ;
 assign um_iw[281] = \col[7].zbuf_top_iw_I[11].z ;
 assign um_iw[282] = \col[7].zbuf_top_iw_I[12].z ;
 assign um_iw[283] = \col[7].zbuf_top_iw_I[13].z ;
 assign um_iw[284] = \col[7].zbuf_top_iw_I[14].z ;
 assign um_iw[285] = \col[7].zbuf_top_iw_I[15].z ;
 assign um_iw[286] = \col[7].zbuf_top_iw_I[16].z ;
 assign um_iw[287] = \col[7].zbuf_top_iw_I[17].z ;
 assign um_iw[271] = \col[7].zbuf_top_iw_I[1].z ;
 assign um_iw[272] = \col[7].zbuf_top_iw_I[2].z ;
 assign um_iw[273] = \col[7].zbuf_top_iw_I[3].z ;
 assign um_iw[274] = \col[7].zbuf_top_iw_I[4].z ;
 assign um_iw[275] = \col[7].zbuf_top_iw_I[5].z ;
 assign um_iw[276] = \col[7].zbuf_top_iw_I[6].z ;
 assign um_iw[277] = \col[7].zbuf_top_iw_I[7].z ;
 assign um_iw[278] = \col[7].zbuf_top_iw_I[8].z ;
 assign um_iw[279] = \col[7].zbuf_top_iw_I[9].z ;
 assign spine_ow[1] = \tbuf_spine_ow_I[0].z ;
 assign spine_ow[11] = \tbuf_spine_ow_I[10].z ;
 assign spine_ow[12] = \tbuf_spine_ow_I[11].z ;
 assign spine_ow[13] = \tbuf_spine_ow_I[12].z ;
 assign spine_ow[14] = \tbuf_spine_ow_I[13].z ;
 assign spine_ow[15] = \tbuf_spine_ow_I[14].z ;
 assign spine_ow[16] = \tbuf_spine_ow_I[15].z ;
 assign spine_ow[17] = \tbuf_spine_ow_I[16].z ;
 assign spine_ow[18] = \tbuf_spine_ow_I[17].z ;
 assign spine_ow[19] = \tbuf_spine_ow_I[18].z ;
 assign spine_ow[20] = \tbuf_spine_ow_I[19].z ;
 assign spine_ow[2] = \tbuf_spine_ow_I[1].z ;
 assign spine_ow[21] = \tbuf_spine_ow_I[20].z ;
 assign spine_ow[22] = \tbuf_spine_ow_I[21].z ;
 assign spine_ow[23] = \tbuf_spine_ow_I[22].z ;
 assign spine_ow[24] = \tbuf_spine_ow_I[23].z ;
 assign spine_ow[3] = \tbuf_spine_ow_I[2].z ;
 assign spine_ow[4] = \tbuf_spine_ow_I[3].z ;
 assign spine_ow[5] = \tbuf_spine_ow_I[4].z ;
 assign spine_ow[6] = \tbuf_spine_ow_I[5].z ;
 assign spine_ow[7] = \tbuf_spine_ow_I[6].z ;
 assign spine_ow[8] = \tbuf_spine_ow_I[7].z ;
 assign spine_ow[9] = \tbuf_spine_ow_I[8].z ;
 assign spine_ow[10] = \tbuf_spine_ow_I[9].z ;
 assign spine_ow[0] = \tie_spine_guard_I[0].lo ;
 assign spine_ow[25] = \tie_spine_guard_I[1].lo ;
endmodule
