module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[1].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[2].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[3].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[4].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[5].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[6].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[0] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[1] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[2] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[3] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[4] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[5] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[6] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uio_out[7] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[0] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[1] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[2] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[3] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[4] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[5] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[6] ;
 wire \top_I.branch[0].col_um[7].um_bot_I.uo_out[7] ;
 wire \top_I.branch[0].l_k_one ;
 wire \top_I.branch[0].l_k_zero ;
 wire \top_I.branch[0].l_um_ena[0] ;
 wire \top_I.branch[0].l_um_ena[10] ;
 wire \top_I.branch[0].l_um_ena[11] ;
 wire \top_I.branch[0].l_um_ena[12] ;
 wire \top_I.branch[0].l_um_ena[13] ;
 wire \top_I.branch[0].l_um_ena[14] ;
 wire \top_I.branch[0].l_um_ena[15] ;
 wire \top_I.branch[0].l_um_ena[1] ;
 wire \top_I.branch[0].l_um_ena[2] ;
 wire \top_I.branch[0].l_um_ena[3] ;
 wire \top_I.branch[0].l_um_ena[4] ;
 wire \top_I.branch[0].l_um_ena[5] ;
 wire \top_I.branch[0].l_um_ena[6] ;
 wire \top_I.branch[0].l_um_ena[7] ;
 wire \top_I.branch[0].l_um_ena[8] ;
 wire \top_I.branch[0].l_um_ena[9] ;
 wire \top_I.branch[0].l_um_iw[0] ;
 wire \top_I.branch[0].l_um_iw[100] ;
 wire \top_I.branch[0].l_um_iw[101] ;
 wire \top_I.branch[0].l_um_iw[102] ;
 wire \top_I.branch[0].l_um_iw[103] ;
 wire \top_I.branch[0].l_um_iw[104] ;
 wire \top_I.branch[0].l_um_iw[105] ;
 wire \top_I.branch[0].l_um_iw[106] ;
 wire \top_I.branch[0].l_um_iw[107] ;
 wire \top_I.branch[0].l_um_iw[108] ;
 wire \top_I.branch[0].l_um_iw[109] ;
 wire \top_I.branch[0].l_um_iw[10] ;
 wire \top_I.branch[0].l_um_iw[110] ;
 wire \top_I.branch[0].l_um_iw[111] ;
 wire \top_I.branch[0].l_um_iw[112] ;
 wire \top_I.branch[0].l_um_iw[113] ;
 wire \top_I.branch[0].l_um_iw[114] ;
 wire \top_I.branch[0].l_um_iw[115] ;
 wire \top_I.branch[0].l_um_iw[116] ;
 wire \top_I.branch[0].l_um_iw[117] ;
 wire \top_I.branch[0].l_um_iw[118] ;
 wire \top_I.branch[0].l_um_iw[119] ;
 wire \top_I.branch[0].l_um_iw[11] ;
 wire \top_I.branch[0].l_um_iw[120] ;
 wire \top_I.branch[0].l_um_iw[121] ;
 wire \top_I.branch[0].l_um_iw[122] ;
 wire \top_I.branch[0].l_um_iw[123] ;
 wire \top_I.branch[0].l_um_iw[124] ;
 wire \top_I.branch[0].l_um_iw[125] ;
 wire \top_I.branch[0].l_um_iw[126] ;
 wire \top_I.branch[0].l_um_iw[127] ;
 wire \top_I.branch[0].l_um_iw[128] ;
 wire \top_I.branch[0].l_um_iw[129] ;
 wire \top_I.branch[0].l_um_iw[12] ;
 wire \top_I.branch[0].l_um_iw[130] ;
 wire \top_I.branch[0].l_um_iw[131] ;
 wire \top_I.branch[0].l_um_iw[132] ;
 wire \top_I.branch[0].l_um_iw[133] ;
 wire \top_I.branch[0].l_um_iw[134] ;
 wire \top_I.branch[0].l_um_iw[135] ;
 wire \top_I.branch[0].l_um_iw[136] ;
 wire \top_I.branch[0].l_um_iw[137] ;
 wire \top_I.branch[0].l_um_iw[138] ;
 wire \top_I.branch[0].l_um_iw[139] ;
 wire \top_I.branch[0].l_um_iw[13] ;
 wire \top_I.branch[0].l_um_iw[140] ;
 wire \top_I.branch[0].l_um_iw[141] ;
 wire \top_I.branch[0].l_um_iw[142] ;
 wire \top_I.branch[0].l_um_iw[143] ;
 wire \top_I.branch[0].l_um_iw[144] ;
 wire \top_I.branch[0].l_um_iw[145] ;
 wire \top_I.branch[0].l_um_iw[146] ;
 wire \top_I.branch[0].l_um_iw[147] ;
 wire \top_I.branch[0].l_um_iw[148] ;
 wire \top_I.branch[0].l_um_iw[149] ;
 wire \top_I.branch[0].l_um_iw[14] ;
 wire \top_I.branch[0].l_um_iw[150] ;
 wire \top_I.branch[0].l_um_iw[151] ;
 wire \top_I.branch[0].l_um_iw[152] ;
 wire \top_I.branch[0].l_um_iw[153] ;
 wire \top_I.branch[0].l_um_iw[154] ;
 wire \top_I.branch[0].l_um_iw[155] ;
 wire \top_I.branch[0].l_um_iw[156] ;
 wire \top_I.branch[0].l_um_iw[157] ;
 wire \top_I.branch[0].l_um_iw[158] ;
 wire \top_I.branch[0].l_um_iw[159] ;
 wire \top_I.branch[0].l_um_iw[15] ;
 wire \top_I.branch[0].l_um_iw[160] ;
 wire \top_I.branch[0].l_um_iw[161] ;
 wire \top_I.branch[0].l_um_iw[162] ;
 wire \top_I.branch[0].l_um_iw[163] ;
 wire \top_I.branch[0].l_um_iw[164] ;
 wire \top_I.branch[0].l_um_iw[165] ;
 wire \top_I.branch[0].l_um_iw[166] ;
 wire \top_I.branch[0].l_um_iw[167] ;
 wire \top_I.branch[0].l_um_iw[168] ;
 wire \top_I.branch[0].l_um_iw[169] ;
 wire \top_I.branch[0].l_um_iw[16] ;
 wire \top_I.branch[0].l_um_iw[170] ;
 wire \top_I.branch[0].l_um_iw[171] ;
 wire \top_I.branch[0].l_um_iw[172] ;
 wire \top_I.branch[0].l_um_iw[173] ;
 wire \top_I.branch[0].l_um_iw[174] ;
 wire \top_I.branch[0].l_um_iw[175] ;
 wire \top_I.branch[0].l_um_iw[176] ;
 wire \top_I.branch[0].l_um_iw[177] ;
 wire \top_I.branch[0].l_um_iw[178] ;
 wire \top_I.branch[0].l_um_iw[179] ;
 wire \top_I.branch[0].l_um_iw[17] ;
 wire \top_I.branch[0].l_um_iw[180] ;
 wire \top_I.branch[0].l_um_iw[181] ;
 wire \top_I.branch[0].l_um_iw[182] ;
 wire \top_I.branch[0].l_um_iw[183] ;
 wire \top_I.branch[0].l_um_iw[184] ;
 wire \top_I.branch[0].l_um_iw[185] ;
 wire \top_I.branch[0].l_um_iw[186] ;
 wire \top_I.branch[0].l_um_iw[187] ;
 wire \top_I.branch[0].l_um_iw[188] ;
 wire \top_I.branch[0].l_um_iw[189] ;
 wire \top_I.branch[0].l_um_iw[18] ;
 wire \top_I.branch[0].l_um_iw[190] ;
 wire \top_I.branch[0].l_um_iw[191] ;
 wire \top_I.branch[0].l_um_iw[192] ;
 wire \top_I.branch[0].l_um_iw[193] ;
 wire \top_I.branch[0].l_um_iw[194] ;
 wire \top_I.branch[0].l_um_iw[195] ;
 wire \top_I.branch[0].l_um_iw[196] ;
 wire \top_I.branch[0].l_um_iw[197] ;
 wire \top_I.branch[0].l_um_iw[198] ;
 wire \top_I.branch[0].l_um_iw[199] ;
 wire \top_I.branch[0].l_um_iw[19] ;
 wire \top_I.branch[0].l_um_iw[1] ;
 wire \top_I.branch[0].l_um_iw[200] ;
 wire \top_I.branch[0].l_um_iw[201] ;
 wire \top_I.branch[0].l_um_iw[202] ;
 wire \top_I.branch[0].l_um_iw[203] ;
 wire \top_I.branch[0].l_um_iw[204] ;
 wire \top_I.branch[0].l_um_iw[205] ;
 wire \top_I.branch[0].l_um_iw[206] ;
 wire \top_I.branch[0].l_um_iw[207] ;
 wire \top_I.branch[0].l_um_iw[208] ;
 wire \top_I.branch[0].l_um_iw[209] ;
 wire \top_I.branch[0].l_um_iw[20] ;
 wire \top_I.branch[0].l_um_iw[210] ;
 wire \top_I.branch[0].l_um_iw[211] ;
 wire \top_I.branch[0].l_um_iw[212] ;
 wire \top_I.branch[0].l_um_iw[213] ;
 wire \top_I.branch[0].l_um_iw[214] ;
 wire \top_I.branch[0].l_um_iw[215] ;
 wire \top_I.branch[0].l_um_iw[216] ;
 wire \top_I.branch[0].l_um_iw[217] ;
 wire \top_I.branch[0].l_um_iw[218] ;
 wire \top_I.branch[0].l_um_iw[219] ;
 wire \top_I.branch[0].l_um_iw[21] ;
 wire \top_I.branch[0].l_um_iw[220] ;
 wire \top_I.branch[0].l_um_iw[221] ;
 wire \top_I.branch[0].l_um_iw[222] ;
 wire \top_I.branch[0].l_um_iw[223] ;
 wire \top_I.branch[0].l_um_iw[224] ;
 wire \top_I.branch[0].l_um_iw[225] ;
 wire \top_I.branch[0].l_um_iw[226] ;
 wire \top_I.branch[0].l_um_iw[227] ;
 wire \top_I.branch[0].l_um_iw[228] ;
 wire \top_I.branch[0].l_um_iw[229] ;
 wire \top_I.branch[0].l_um_iw[22] ;
 wire \top_I.branch[0].l_um_iw[230] ;
 wire \top_I.branch[0].l_um_iw[231] ;
 wire \top_I.branch[0].l_um_iw[232] ;
 wire \top_I.branch[0].l_um_iw[233] ;
 wire \top_I.branch[0].l_um_iw[234] ;
 wire \top_I.branch[0].l_um_iw[235] ;
 wire \top_I.branch[0].l_um_iw[236] ;
 wire \top_I.branch[0].l_um_iw[237] ;
 wire \top_I.branch[0].l_um_iw[238] ;
 wire \top_I.branch[0].l_um_iw[239] ;
 wire \top_I.branch[0].l_um_iw[23] ;
 wire \top_I.branch[0].l_um_iw[240] ;
 wire \top_I.branch[0].l_um_iw[241] ;
 wire \top_I.branch[0].l_um_iw[242] ;
 wire \top_I.branch[0].l_um_iw[243] ;
 wire \top_I.branch[0].l_um_iw[244] ;
 wire \top_I.branch[0].l_um_iw[245] ;
 wire \top_I.branch[0].l_um_iw[246] ;
 wire \top_I.branch[0].l_um_iw[247] ;
 wire \top_I.branch[0].l_um_iw[248] ;
 wire \top_I.branch[0].l_um_iw[249] ;
 wire \top_I.branch[0].l_um_iw[24] ;
 wire \top_I.branch[0].l_um_iw[250] ;
 wire \top_I.branch[0].l_um_iw[251] ;
 wire \top_I.branch[0].l_um_iw[252] ;
 wire \top_I.branch[0].l_um_iw[253] ;
 wire \top_I.branch[0].l_um_iw[254] ;
 wire \top_I.branch[0].l_um_iw[255] ;
 wire \top_I.branch[0].l_um_iw[256] ;
 wire \top_I.branch[0].l_um_iw[257] ;
 wire \top_I.branch[0].l_um_iw[258] ;
 wire \top_I.branch[0].l_um_iw[259] ;
 wire \top_I.branch[0].l_um_iw[25] ;
 wire \top_I.branch[0].l_um_iw[260] ;
 wire \top_I.branch[0].l_um_iw[261] ;
 wire \top_I.branch[0].l_um_iw[262] ;
 wire \top_I.branch[0].l_um_iw[263] ;
 wire \top_I.branch[0].l_um_iw[264] ;
 wire \top_I.branch[0].l_um_iw[265] ;
 wire \top_I.branch[0].l_um_iw[266] ;
 wire \top_I.branch[0].l_um_iw[267] ;
 wire \top_I.branch[0].l_um_iw[268] ;
 wire \top_I.branch[0].l_um_iw[269] ;
 wire \top_I.branch[0].l_um_iw[26] ;
 wire \top_I.branch[0].l_um_iw[270] ;
 wire \top_I.branch[0].l_um_iw[271] ;
 wire \top_I.branch[0].l_um_iw[272] ;
 wire \top_I.branch[0].l_um_iw[273] ;
 wire \top_I.branch[0].l_um_iw[274] ;
 wire \top_I.branch[0].l_um_iw[275] ;
 wire \top_I.branch[0].l_um_iw[276] ;
 wire \top_I.branch[0].l_um_iw[277] ;
 wire \top_I.branch[0].l_um_iw[278] ;
 wire \top_I.branch[0].l_um_iw[279] ;
 wire \top_I.branch[0].l_um_iw[27] ;
 wire \top_I.branch[0].l_um_iw[280] ;
 wire \top_I.branch[0].l_um_iw[281] ;
 wire \top_I.branch[0].l_um_iw[282] ;
 wire \top_I.branch[0].l_um_iw[283] ;
 wire \top_I.branch[0].l_um_iw[284] ;
 wire \top_I.branch[0].l_um_iw[285] ;
 wire \top_I.branch[0].l_um_iw[286] ;
 wire \top_I.branch[0].l_um_iw[287] ;
 wire \top_I.branch[0].l_um_iw[28] ;
 wire \top_I.branch[0].l_um_iw[29] ;
 wire \top_I.branch[0].l_um_iw[2] ;
 wire \top_I.branch[0].l_um_iw[30] ;
 wire \top_I.branch[0].l_um_iw[31] ;
 wire \top_I.branch[0].l_um_iw[32] ;
 wire \top_I.branch[0].l_um_iw[33] ;
 wire \top_I.branch[0].l_um_iw[34] ;
 wire \top_I.branch[0].l_um_iw[35] ;
 wire \top_I.branch[0].l_um_iw[36] ;
 wire \top_I.branch[0].l_um_iw[37] ;
 wire \top_I.branch[0].l_um_iw[38] ;
 wire \top_I.branch[0].l_um_iw[39] ;
 wire \top_I.branch[0].l_um_iw[3] ;
 wire \top_I.branch[0].l_um_iw[40] ;
 wire \top_I.branch[0].l_um_iw[41] ;
 wire \top_I.branch[0].l_um_iw[42] ;
 wire \top_I.branch[0].l_um_iw[43] ;
 wire \top_I.branch[0].l_um_iw[44] ;
 wire \top_I.branch[0].l_um_iw[45] ;
 wire \top_I.branch[0].l_um_iw[46] ;
 wire \top_I.branch[0].l_um_iw[47] ;
 wire \top_I.branch[0].l_um_iw[48] ;
 wire \top_I.branch[0].l_um_iw[49] ;
 wire \top_I.branch[0].l_um_iw[4] ;
 wire \top_I.branch[0].l_um_iw[50] ;
 wire \top_I.branch[0].l_um_iw[51] ;
 wire \top_I.branch[0].l_um_iw[52] ;
 wire \top_I.branch[0].l_um_iw[53] ;
 wire \top_I.branch[0].l_um_iw[54] ;
 wire \top_I.branch[0].l_um_iw[55] ;
 wire \top_I.branch[0].l_um_iw[56] ;
 wire \top_I.branch[0].l_um_iw[57] ;
 wire \top_I.branch[0].l_um_iw[58] ;
 wire \top_I.branch[0].l_um_iw[59] ;
 wire \top_I.branch[0].l_um_iw[5] ;
 wire \top_I.branch[0].l_um_iw[60] ;
 wire \top_I.branch[0].l_um_iw[61] ;
 wire \top_I.branch[0].l_um_iw[62] ;
 wire \top_I.branch[0].l_um_iw[63] ;
 wire \top_I.branch[0].l_um_iw[64] ;
 wire \top_I.branch[0].l_um_iw[65] ;
 wire \top_I.branch[0].l_um_iw[66] ;
 wire \top_I.branch[0].l_um_iw[67] ;
 wire \top_I.branch[0].l_um_iw[68] ;
 wire \top_I.branch[0].l_um_iw[69] ;
 wire \top_I.branch[0].l_um_iw[6] ;
 wire \top_I.branch[0].l_um_iw[70] ;
 wire \top_I.branch[0].l_um_iw[71] ;
 wire \top_I.branch[0].l_um_iw[72] ;
 wire \top_I.branch[0].l_um_iw[73] ;
 wire \top_I.branch[0].l_um_iw[74] ;
 wire \top_I.branch[0].l_um_iw[75] ;
 wire \top_I.branch[0].l_um_iw[76] ;
 wire \top_I.branch[0].l_um_iw[77] ;
 wire \top_I.branch[0].l_um_iw[78] ;
 wire \top_I.branch[0].l_um_iw[79] ;
 wire \top_I.branch[0].l_um_iw[7] ;
 wire \top_I.branch[0].l_um_iw[80] ;
 wire \top_I.branch[0].l_um_iw[81] ;
 wire \top_I.branch[0].l_um_iw[82] ;
 wire \top_I.branch[0].l_um_iw[83] ;
 wire \top_I.branch[0].l_um_iw[84] ;
 wire \top_I.branch[0].l_um_iw[85] ;
 wire \top_I.branch[0].l_um_iw[86] ;
 wire \top_I.branch[0].l_um_iw[87] ;
 wire \top_I.branch[0].l_um_iw[88] ;
 wire \top_I.branch[0].l_um_iw[89] ;
 wire \top_I.branch[0].l_um_iw[8] ;
 wire \top_I.branch[0].l_um_iw[90] ;
 wire \top_I.branch[0].l_um_iw[91] ;
 wire \top_I.branch[0].l_um_iw[92] ;
 wire \top_I.branch[0].l_um_iw[93] ;
 wire \top_I.branch[0].l_um_iw[94] ;
 wire \top_I.branch[0].l_um_iw[95] ;
 wire \top_I.branch[0].l_um_iw[96] ;
 wire \top_I.branch[0].l_um_iw[97] ;
 wire \top_I.branch[0].l_um_iw[98] ;
 wire \top_I.branch[0].l_um_iw[99] ;
 wire \top_I.branch[0].l_um_iw[9] ;
 wire \top_I.branch[0].l_um_k_zero[0] ;
 wire \top_I.branch[0].l_um_k_zero[10] ;
 wire \top_I.branch[0].l_um_k_zero[11] ;
 wire \top_I.branch[0].l_um_k_zero[12] ;
 wire \top_I.branch[0].l_um_k_zero[13] ;
 wire \top_I.branch[0].l_um_k_zero[14] ;
 wire \top_I.branch[0].l_um_k_zero[15] ;
 wire \top_I.branch[0].l_um_k_zero[1] ;
 wire \top_I.branch[0].l_um_k_zero[2] ;
 wire \top_I.branch[0].l_um_k_zero[3] ;
 wire \top_I.branch[0].l_um_k_zero[4] ;
 wire \top_I.branch[0].l_um_k_zero[5] ;
 wire \top_I.branch[0].l_um_k_zero[6] ;
 wire \top_I.branch[0].l_um_k_zero[7] ;
 wire \top_I.branch[0].l_um_k_zero[8] ;
 wire \top_I.branch[0].l_um_k_zero[9] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[10].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[10].l_k_one ;
 wire \top_I.branch[10].l_k_zero ;
 wire \top_I.branch[10].l_um_ena[0] ;
 wire \top_I.branch[10].l_um_ena[10] ;
 wire \top_I.branch[10].l_um_ena[11] ;
 wire \top_I.branch[10].l_um_ena[12] ;
 wire \top_I.branch[10].l_um_ena[13] ;
 wire \top_I.branch[10].l_um_ena[14] ;
 wire \top_I.branch[10].l_um_ena[15] ;
 wire \top_I.branch[10].l_um_ena[1] ;
 wire \top_I.branch[10].l_um_ena[2] ;
 wire \top_I.branch[10].l_um_ena[3] ;
 wire \top_I.branch[10].l_um_ena[4] ;
 wire \top_I.branch[10].l_um_ena[5] ;
 wire \top_I.branch[10].l_um_ena[6] ;
 wire \top_I.branch[10].l_um_ena[7] ;
 wire \top_I.branch[10].l_um_ena[8] ;
 wire \top_I.branch[10].l_um_ena[9] ;
 wire \top_I.branch[10].l_um_iw[0] ;
 wire \top_I.branch[10].l_um_iw[100] ;
 wire \top_I.branch[10].l_um_iw[101] ;
 wire \top_I.branch[10].l_um_iw[102] ;
 wire \top_I.branch[10].l_um_iw[103] ;
 wire \top_I.branch[10].l_um_iw[104] ;
 wire \top_I.branch[10].l_um_iw[105] ;
 wire \top_I.branch[10].l_um_iw[106] ;
 wire \top_I.branch[10].l_um_iw[107] ;
 wire \top_I.branch[10].l_um_iw[108] ;
 wire \top_I.branch[10].l_um_iw[109] ;
 wire \top_I.branch[10].l_um_iw[10] ;
 wire \top_I.branch[10].l_um_iw[110] ;
 wire \top_I.branch[10].l_um_iw[111] ;
 wire \top_I.branch[10].l_um_iw[112] ;
 wire \top_I.branch[10].l_um_iw[113] ;
 wire \top_I.branch[10].l_um_iw[114] ;
 wire \top_I.branch[10].l_um_iw[115] ;
 wire \top_I.branch[10].l_um_iw[116] ;
 wire \top_I.branch[10].l_um_iw[117] ;
 wire \top_I.branch[10].l_um_iw[118] ;
 wire \top_I.branch[10].l_um_iw[119] ;
 wire \top_I.branch[10].l_um_iw[11] ;
 wire \top_I.branch[10].l_um_iw[120] ;
 wire \top_I.branch[10].l_um_iw[121] ;
 wire \top_I.branch[10].l_um_iw[122] ;
 wire \top_I.branch[10].l_um_iw[123] ;
 wire \top_I.branch[10].l_um_iw[124] ;
 wire \top_I.branch[10].l_um_iw[125] ;
 wire \top_I.branch[10].l_um_iw[126] ;
 wire \top_I.branch[10].l_um_iw[127] ;
 wire \top_I.branch[10].l_um_iw[128] ;
 wire \top_I.branch[10].l_um_iw[129] ;
 wire \top_I.branch[10].l_um_iw[12] ;
 wire \top_I.branch[10].l_um_iw[130] ;
 wire \top_I.branch[10].l_um_iw[131] ;
 wire \top_I.branch[10].l_um_iw[132] ;
 wire \top_I.branch[10].l_um_iw[133] ;
 wire \top_I.branch[10].l_um_iw[134] ;
 wire \top_I.branch[10].l_um_iw[135] ;
 wire \top_I.branch[10].l_um_iw[136] ;
 wire \top_I.branch[10].l_um_iw[137] ;
 wire \top_I.branch[10].l_um_iw[138] ;
 wire \top_I.branch[10].l_um_iw[139] ;
 wire \top_I.branch[10].l_um_iw[13] ;
 wire \top_I.branch[10].l_um_iw[140] ;
 wire \top_I.branch[10].l_um_iw[141] ;
 wire \top_I.branch[10].l_um_iw[142] ;
 wire \top_I.branch[10].l_um_iw[143] ;
 wire \top_I.branch[10].l_um_iw[144] ;
 wire \top_I.branch[10].l_um_iw[145] ;
 wire \top_I.branch[10].l_um_iw[146] ;
 wire \top_I.branch[10].l_um_iw[147] ;
 wire \top_I.branch[10].l_um_iw[148] ;
 wire \top_I.branch[10].l_um_iw[149] ;
 wire \top_I.branch[10].l_um_iw[14] ;
 wire \top_I.branch[10].l_um_iw[150] ;
 wire \top_I.branch[10].l_um_iw[151] ;
 wire \top_I.branch[10].l_um_iw[152] ;
 wire \top_I.branch[10].l_um_iw[153] ;
 wire \top_I.branch[10].l_um_iw[154] ;
 wire \top_I.branch[10].l_um_iw[155] ;
 wire \top_I.branch[10].l_um_iw[156] ;
 wire \top_I.branch[10].l_um_iw[157] ;
 wire \top_I.branch[10].l_um_iw[158] ;
 wire \top_I.branch[10].l_um_iw[159] ;
 wire \top_I.branch[10].l_um_iw[15] ;
 wire \top_I.branch[10].l_um_iw[160] ;
 wire \top_I.branch[10].l_um_iw[161] ;
 wire \top_I.branch[10].l_um_iw[162] ;
 wire \top_I.branch[10].l_um_iw[163] ;
 wire \top_I.branch[10].l_um_iw[164] ;
 wire \top_I.branch[10].l_um_iw[165] ;
 wire \top_I.branch[10].l_um_iw[166] ;
 wire \top_I.branch[10].l_um_iw[167] ;
 wire \top_I.branch[10].l_um_iw[168] ;
 wire \top_I.branch[10].l_um_iw[169] ;
 wire \top_I.branch[10].l_um_iw[16] ;
 wire \top_I.branch[10].l_um_iw[170] ;
 wire \top_I.branch[10].l_um_iw[171] ;
 wire \top_I.branch[10].l_um_iw[172] ;
 wire \top_I.branch[10].l_um_iw[173] ;
 wire \top_I.branch[10].l_um_iw[174] ;
 wire \top_I.branch[10].l_um_iw[175] ;
 wire \top_I.branch[10].l_um_iw[176] ;
 wire \top_I.branch[10].l_um_iw[177] ;
 wire \top_I.branch[10].l_um_iw[178] ;
 wire \top_I.branch[10].l_um_iw[179] ;
 wire \top_I.branch[10].l_um_iw[17] ;
 wire \top_I.branch[10].l_um_iw[180] ;
 wire \top_I.branch[10].l_um_iw[181] ;
 wire \top_I.branch[10].l_um_iw[182] ;
 wire \top_I.branch[10].l_um_iw[183] ;
 wire \top_I.branch[10].l_um_iw[184] ;
 wire \top_I.branch[10].l_um_iw[185] ;
 wire \top_I.branch[10].l_um_iw[186] ;
 wire \top_I.branch[10].l_um_iw[187] ;
 wire \top_I.branch[10].l_um_iw[188] ;
 wire \top_I.branch[10].l_um_iw[189] ;
 wire \top_I.branch[10].l_um_iw[18] ;
 wire \top_I.branch[10].l_um_iw[190] ;
 wire \top_I.branch[10].l_um_iw[191] ;
 wire \top_I.branch[10].l_um_iw[192] ;
 wire \top_I.branch[10].l_um_iw[193] ;
 wire \top_I.branch[10].l_um_iw[194] ;
 wire \top_I.branch[10].l_um_iw[195] ;
 wire \top_I.branch[10].l_um_iw[196] ;
 wire \top_I.branch[10].l_um_iw[197] ;
 wire \top_I.branch[10].l_um_iw[198] ;
 wire \top_I.branch[10].l_um_iw[199] ;
 wire \top_I.branch[10].l_um_iw[19] ;
 wire \top_I.branch[10].l_um_iw[1] ;
 wire \top_I.branch[10].l_um_iw[200] ;
 wire \top_I.branch[10].l_um_iw[201] ;
 wire \top_I.branch[10].l_um_iw[202] ;
 wire \top_I.branch[10].l_um_iw[203] ;
 wire \top_I.branch[10].l_um_iw[204] ;
 wire \top_I.branch[10].l_um_iw[205] ;
 wire \top_I.branch[10].l_um_iw[206] ;
 wire \top_I.branch[10].l_um_iw[207] ;
 wire \top_I.branch[10].l_um_iw[208] ;
 wire \top_I.branch[10].l_um_iw[209] ;
 wire \top_I.branch[10].l_um_iw[20] ;
 wire \top_I.branch[10].l_um_iw[210] ;
 wire \top_I.branch[10].l_um_iw[211] ;
 wire \top_I.branch[10].l_um_iw[212] ;
 wire \top_I.branch[10].l_um_iw[213] ;
 wire \top_I.branch[10].l_um_iw[214] ;
 wire \top_I.branch[10].l_um_iw[215] ;
 wire \top_I.branch[10].l_um_iw[216] ;
 wire \top_I.branch[10].l_um_iw[217] ;
 wire \top_I.branch[10].l_um_iw[218] ;
 wire \top_I.branch[10].l_um_iw[219] ;
 wire \top_I.branch[10].l_um_iw[21] ;
 wire \top_I.branch[10].l_um_iw[220] ;
 wire \top_I.branch[10].l_um_iw[221] ;
 wire \top_I.branch[10].l_um_iw[222] ;
 wire \top_I.branch[10].l_um_iw[223] ;
 wire \top_I.branch[10].l_um_iw[224] ;
 wire \top_I.branch[10].l_um_iw[225] ;
 wire \top_I.branch[10].l_um_iw[226] ;
 wire \top_I.branch[10].l_um_iw[227] ;
 wire \top_I.branch[10].l_um_iw[228] ;
 wire \top_I.branch[10].l_um_iw[229] ;
 wire \top_I.branch[10].l_um_iw[22] ;
 wire \top_I.branch[10].l_um_iw[230] ;
 wire \top_I.branch[10].l_um_iw[231] ;
 wire \top_I.branch[10].l_um_iw[232] ;
 wire \top_I.branch[10].l_um_iw[233] ;
 wire \top_I.branch[10].l_um_iw[234] ;
 wire \top_I.branch[10].l_um_iw[235] ;
 wire \top_I.branch[10].l_um_iw[236] ;
 wire \top_I.branch[10].l_um_iw[237] ;
 wire \top_I.branch[10].l_um_iw[238] ;
 wire \top_I.branch[10].l_um_iw[239] ;
 wire \top_I.branch[10].l_um_iw[23] ;
 wire \top_I.branch[10].l_um_iw[240] ;
 wire \top_I.branch[10].l_um_iw[241] ;
 wire \top_I.branch[10].l_um_iw[242] ;
 wire \top_I.branch[10].l_um_iw[243] ;
 wire \top_I.branch[10].l_um_iw[244] ;
 wire \top_I.branch[10].l_um_iw[245] ;
 wire \top_I.branch[10].l_um_iw[246] ;
 wire \top_I.branch[10].l_um_iw[247] ;
 wire \top_I.branch[10].l_um_iw[248] ;
 wire \top_I.branch[10].l_um_iw[249] ;
 wire \top_I.branch[10].l_um_iw[24] ;
 wire \top_I.branch[10].l_um_iw[250] ;
 wire \top_I.branch[10].l_um_iw[251] ;
 wire \top_I.branch[10].l_um_iw[252] ;
 wire \top_I.branch[10].l_um_iw[253] ;
 wire \top_I.branch[10].l_um_iw[254] ;
 wire \top_I.branch[10].l_um_iw[255] ;
 wire \top_I.branch[10].l_um_iw[256] ;
 wire \top_I.branch[10].l_um_iw[257] ;
 wire \top_I.branch[10].l_um_iw[258] ;
 wire \top_I.branch[10].l_um_iw[259] ;
 wire \top_I.branch[10].l_um_iw[25] ;
 wire \top_I.branch[10].l_um_iw[260] ;
 wire \top_I.branch[10].l_um_iw[261] ;
 wire \top_I.branch[10].l_um_iw[262] ;
 wire \top_I.branch[10].l_um_iw[263] ;
 wire \top_I.branch[10].l_um_iw[264] ;
 wire \top_I.branch[10].l_um_iw[265] ;
 wire \top_I.branch[10].l_um_iw[266] ;
 wire \top_I.branch[10].l_um_iw[267] ;
 wire \top_I.branch[10].l_um_iw[268] ;
 wire \top_I.branch[10].l_um_iw[269] ;
 wire \top_I.branch[10].l_um_iw[26] ;
 wire \top_I.branch[10].l_um_iw[270] ;
 wire \top_I.branch[10].l_um_iw[271] ;
 wire \top_I.branch[10].l_um_iw[272] ;
 wire \top_I.branch[10].l_um_iw[273] ;
 wire \top_I.branch[10].l_um_iw[274] ;
 wire \top_I.branch[10].l_um_iw[275] ;
 wire \top_I.branch[10].l_um_iw[276] ;
 wire \top_I.branch[10].l_um_iw[277] ;
 wire \top_I.branch[10].l_um_iw[278] ;
 wire \top_I.branch[10].l_um_iw[279] ;
 wire \top_I.branch[10].l_um_iw[27] ;
 wire \top_I.branch[10].l_um_iw[280] ;
 wire \top_I.branch[10].l_um_iw[281] ;
 wire \top_I.branch[10].l_um_iw[282] ;
 wire \top_I.branch[10].l_um_iw[283] ;
 wire \top_I.branch[10].l_um_iw[284] ;
 wire \top_I.branch[10].l_um_iw[285] ;
 wire \top_I.branch[10].l_um_iw[286] ;
 wire \top_I.branch[10].l_um_iw[287] ;
 wire \top_I.branch[10].l_um_iw[28] ;
 wire \top_I.branch[10].l_um_iw[29] ;
 wire \top_I.branch[10].l_um_iw[2] ;
 wire \top_I.branch[10].l_um_iw[30] ;
 wire \top_I.branch[10].l_um_iw[31] ;
 wire \top_I.branch[10].l_um_iw[32] ;
 wire \top_I.branch[10].l_um_iw[33] ;
 wire \top_I.branch[10].l_um_iw[34] ;
 wire \top_I.branch[10].l_um_iw[35] ;
 wire \top_I.branch[10].l_um_iw[36] ;
 wire \top_I.branch[10].l_um_iw[37] ;
 wire \top_I.branch[10].l_um_iw[38] ;
 wire \top_I.branch[10].l_um_iw[39] ;
 wire \top_I.branch[10].l_um_iw[3] ;
 wire \top_I.branch[10].l_um_iw[40] ;
 wire \top_I.branch[10].l_um_iw[41] ;
 wire \top_I.branch[10].l_um_iw[42] ;
 wire \top_I.branch[10].l_um_iw[43] ;
 wire \top_I.branch[10].l_um_iw[44] ;
 wire \top_I.branch[10].l_um_iw[45] ;
 wire \top_I.branch[10].l_um_iw[46] ;
 wire \top_I.branch[10].l_um_iw[47] ;
 wire \top_I.branch[10].l_um_iw[48] ;
 wire \top_I.branch[10].l_um_iw[49] ;
 wire \top_I.branch[10].l_um_iw[4] ;
 wire \top_I.branch[10].l_um_iw[50] ;
 wire \top_I.branch[10].l_um_iw[51] ;
 wire \top_I.branch[10].l_um_iw[52] ;
 wire \top_I.branch[10].l_um_iw[53] ;
 wire \top_I.branch[10].l_um_iw[54] ;
 wire \top_I.branch[10].l_um_iw[55] ;
 wire \top_I.branch[10].l_um_iw[56] ;
 wire \top_I.branch[10].l_um_iw[57] ;
 wire \top_I.branch[10].l_um_iw[58] ;
 wire \top_I.branch[10].l_um_iw[59] ;
 wire \top_I.branch[10].l_um_iw[5] ;
 wire \top_I.branch[10].l_um_iw[60] ;
 wire \top_I.branch[10].l_um_iw[61] ;
 wire \top_I.branch[10].l_um_iw[62] ;
 wire \top_I.branch[10].l_um_iw[63] ;
 wire \top_I.branch[10].l_um_iw[64] ;
 wire \top_I.branch[10].l_um_iw[65] ;
 wire \top_I.branch[10].l_um_iw[66] ;
 wire \top_I.branch[10].l_um_iw[67] ;
 wire \top_I.branch[10].l_um_iw[68] ;
 wire \top_I.branch[10].l_um_iw[69] ;
 wire \top_I.branch[10].l_um_iw[6] ;
 wire \top_I.branch[10].l_um_iw[70] ;
 wire \top_I.branch[10].l_um_iw[71] ;
 wire \top_I.branch[10].l_um_iw[72] ;
 wire \top_I.branch[10].l_um_iw[73] ;
 wire \top_I.branch[10].l_um_iw[74] ;
 wire \top_I.branch[10].l_um_iw[75] ;
 wire \top_I.branch[10].l_um_iw[76] ;
 wire \top_I.branch[10].l_um_iw[77] ;
 wire \top_I.branch[10].l_um_iw[78] ;
 wire \top_I.branch[10].l_um_iw[79] ;
 wire \top_I.branch[10].l_um_iw[7] ;
 wire \top_I.branch[10].l_um_iw[80] ;
 wire \top_I.branch[10].l_um_iw[81] ;
 wire \top_I.branch[10].l_um_iw[82] ;
 wire \top_I.branch[10].l_um_iw[83] ;
 wire \top_I.branch[10].l_um_iw[84] ;
 wire \top_I.branch[10].l_um_iw[85] ;
 wire \top_I.branch[10].l_um_iw[86] ;
 wire \top_I.branch[10].l_um_iw[87] ;
 wire \top_I.branch[10].l_um_iw[88] ;
 wire \top_I.branch[10].l_um_iw[89] ;
 wire \top_I.branch[10].l_um_iw[8] ;
 wire \top_I.branch[10].l_um_iw[90] ;
 wire \top_I.branch[10].l_um_iw[91] ;
 wire \top_I.branch[10].l_um_iw[92] ;
 wire \top_I.branch[10].l_um_iw[93] ;
 wire \top_I.branch[10].l_um_iw[94] ;
 wire \top_I.branch[10].l_um_iw[95] ;
 wire \top_I.branch[10].l_um_iw[96] ;
 wire \top_I.branch[10].l_um_iw[97] ;
 wire \top_I.branch[10].l_um_iw[98] ;
 wire \top_I.branch[10].l_um_iw[99] ;
 wire \top_I.branch[10].l_um_iw[9] ;
 wire \top_I.branch[10].l_um_k_zero[0] ;
 wire \top_I.branch[10].l_um_k_zero[10] ;
 wire \top_I.branch[10].l_um_k_zero[11] ;
 wire \top_I.branch[10].l_um_k_zero[12] ;
 wire \top_I.branch[10].l_um_k_zero[13] ;
 wire \top_I.branch[10].l_um_k_zero[14] ;
 wire \top_I.branch[10].l_um_k_zero[15] ;
 wire \top_I.branch[10].l_um_k_zero[1] ;
 wire \top_I.branch[10].l_um_k_zero[2] ;
 wire \top_I.branch[10].l_um_k_zero[3] ;
 wire \top_I.branch[10].l_um_k_zero[4] ;
 wire \top_I.branch[10].l_um_k_zero[5] ;
 wire \top_I.branch[10].l_um_k_zero[6] ;
 wire \top_I.branch[10].l_um_k_zero[7] ;
 wire \top_I.branch[10].l_um_k_zero[8] ;
 wire \top_I.branch[10].l_um_k_zero[9] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[11].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[11].l_k_one ;
 wire \top_I.branch[11].l_k_zero ;
 wire \top_I.branch[11].l_um_ena[0] ;
 wire \top_I.branch[11].l_um_ena[10] ;
 wire \top_I.branch[11].l_um_ena[11] ;
 wire \top_I.branch[11].l_um_ena[12] ;
 wire \top_I.branch[11].l_um_ena[13] ;
 wire \top_I.branch[11].l_um_ena[14] ;
 wire \top_I.branch[11].l_um_ena[15] ;
 wire \top_I.branch[11].l_um_ena[1] ;
 wire \top_I.branch[11].l_um_ena[2] ;
 wire \top_I.branch[11].l_um_ena[3] ;
 wire \top_I.branch[11].l_um_ena[4] ;
 wire \top_I.branch[11].l_um_ena[5] ;
 wire \top_I.branch[11].l_um_ena[6] ;
 wire \top_I.branch[11].l_um_ena[7] ;
 wire \top_I.branch[11].l_um_ena[8] ;
 wire \top_I.branch[11].l_um_ena[9] ;
 wire \top_I.branch[11].l_um_iw[0] ;
 wire \top_I.branch[11].l_um_iw[100] ;
 wire \top_I.branch[11].l_um_iw[101] ;
 wire \top_I.branch[11].l_um_iw[102] ;
 wire \top_I.branch[11].l_um_iw[103] ;
 wire \top_I.branch[11].l_um_iw[104] ;
 wire \top_I.branch[11].l_um_iw[105] ;
 wire \top_I.branch[11].l_um_iw[106] ;
 wire \top_I.branch[11].l_um_iw[107] ;
 wire \top_I.branch[11].l_um_iw[108] ;
 wire \top_I.branch[11].l_um_iw[109] ;
 wire \top_I.branch[11].l_um_iw[10] ;
 wire \top_I.branch[11].l_um_iw[110] ;
 wire \top_I.branch[11].l_um_iw[111] ;
 wire \top_I.branch[11].l_um_iw[112] ;
 wire \top_I.branch[11].l_um_iw[113] ;
 wire \top_I.branch[11].l_um_iw[114] ;
 wire \top_I.branch[11].l_um_iw[115] ;
 wire \top_I.branch[11].l_um_iw[116] ;
 wire \top_I.branch[11].l_um_iw[117] ;
 wire \top_I.branch[11].l_um_iw[118] ;
 wire \top_I.branch[11].l_um_iw[119] ;
 wire \top_I.branch[11].l_um_iw[11] ;
 wire \top_I.branch[11].l_um_iw[120] ;
 wire \top_I.branch[11].l_um_iw[121] ;
 wire \top_I.branch[11].l_um_iw[122] ;
 wire \top_I.branch[11].l_um_iw[123] ;
 wire \top_I.branch[11].l_um_iw[124] ;
 wire \top_I.branch[11].l_um_iw[125] ;
 wire \top_I.branch[11].l_um_iw[126] ;
 wire \top_I.branch[11].l_um_iw[127] ;
 wire \top_I.branch[11].l_um_iw[128] ;
 wire \top_I.branch[11].l_um_iw[129] ;
 wire \top_I.branch[11].l_um_iw[12] ;
 wire \top_I.branch[11].l_um_iw[130] ;
 wire \top_I.branch[11].l_um_iw[131] ;
 wire \top_I.branch[11].l_um_iw[132] ;
 wire \top_I.branch[11].l_um_iw[133] ;
 wire \top_I.branch[11].l_um_iw[134] ;
 wire \top_I.branch[11].l_um_iw[135] ;
 wire \top_I.branch[11].l_um_iw[136] ;
 wire \top_I.branch[11].l_um_iw[137] ;
 wire \top_I.branch[11].l_um_iw[138] ;
 wire \top_I.branch[11].l_um_iw[139] ;
 wire \top_I.branch[11].l_um_iw[13] ;
 wire \top_I.branch[11].l_um_iw[140] ;
 wire \top_I.branch[11].l_um_iw[141] ;
 wire \top_I.branch[11].l_um_iw[142] ;
 wire \top_I.branch[11].l_um_iw[143] ;
 wire \top_I.branch[11].l_um_iw[144] ;
 wire \top_I.branch[11].l_um_iw[145] ;
 wire \top_I.branch[11].l_um_iw[146] ;
 wire \top_I.branch[11].l_um_iw[147] ;
 wire \top_I.branch[11].l_um_iw[148] ;
 wire \top_I.branch[11].l_um_iw[149] ;
 wire \top_I.branch[11].l_um_iw[14] ;
 wire \top_I.branch[11].l_um_iw[150] ;
 wire \top_I.branch[11].l_um_iw[151] ;
 wire \top_I.branch[11].l_um_iw[152] ;
 wire \top_I.branch[11].l_um_iw[153] ;
 wire \top_I.branch[11].l_um_iw[154] ;
 wire \top_I.branch[11].l_um_iw[155] ;
 wire \top_I.branch[11].l_um_iw[156] ;
 wire \top_I.branch[11].l_um_iw[157] ;
 wire \top_I.branch[11].l_um_iw[158] ;
 wire \top_I.branch[11].l_um_iw[159] ;
 wire \top_I.branch[11].l_um_iw[15] ;
 wire \top_I.branch[11].l_um_iw[160] ;
 wire \top_I.branch[11].l_um_iw[161] ;
 wire \top_I.branch[11].l_um_iw[162] ;
 wire \top_I.branch[11].l_um_iw[163] ;
 wire \top_I.branch[11].l_um_iw[164] ;
 wire \top_I.branch[11].l_um_iw[165] ;
 wire \top_I.branch[11].l_um_iw[166] ;
 wire \top_I.branch[11].l_um_iw[167] ;
 wire \top_I.branch[11].l_um_iw[168] ;
 wire \top_I.branch[11].l_um_iw[169] ;
 wire \top_I.branch[11].l_um_iw[16] ;
 wire \top_I.branch[11].l_um_iw[170] ;
 wire \top_I.branch[11].l_um_iw[171] ;
 wire \top_I.branch[11].l_um_iw[172] ;
 wire \top_I.branch[11].l_um_iw[173] ;
 wire \top_I.branch[11].l_um_iw[174] ;
 wire \top_I.branch[11].l_um_iw[175] ;
 wire \top_I.branch[11].l_um_iw[176] ;
 wire \top_I.branch[11].l_um_iw[177] ;
 wire \top_I.branch[11].l_um_iw[178] ;
 wire \top_I.branch[11].l_um_iw[179] ;
 wire \top_I.branch[11].l_um_iw[17] ;
 wire \top_I.branch[11].l_um_iw[180] ;
 wire \top_I.branch[11].l_um_iw[181] ;
 wire \top_I.branch[11].l_um_iw[182] ;
 wire \top_I.branch[11].l_um_iw[183] ;
 wire \top_I.branch[11].l_um_iw[184] ;
 wire \top_I.branch[11].l_um_iw[185] ;
 wire \top_I.branch[11].l_um_iw[186] ;
 wire \top_I.branch[11].l_um_iw[187] ;
 wire \top_I.branch[11].l_um_iw[188] ;
 wire \top_I.branch[11].l_um_iw[189] ;
 wire \top_I.branch[11].l_um_iw[18] ;
 wire \top_I.branch[11].l_um_iw[190] ;
 wire \top_I.branch[11].l_um_iw[191] ;
 wire \top_I.branch[11].l_um_iw[192] ;
 wire \top_I.branch[11].l_um_iw[193] ;
 wire \top_I.branch[11].l_um_iw[194] ;
 wire \top_I.branch[11].l_um_iw[195] ;
 wire \top_I.branch[11].l_um_iw[196] ;
 wire \top_I.branch[11].l_um_iw[197] ;
 wire \top_I.branch[11].l_um_iw[198] ;
 wire \top_I.branch[11].l_um_iw[199] ;
 wire \top_I.branch[11].l_um_iw[19] ;
 wire \top_I.branch[11].l_um_iw[1] ;
 wire \top_I.branch[11].l_um_iw[200] ;
 wire \top_I.branch[11].l_um_iw[201] ;
 wire \top_I.branch[11].l_um_iw[202] ;
 wire \top_I.branch[11].l_um_iw[203] ;
 wire \top_I.branch[11].l_um_iw[204] ;
 wire \top_I.branch[11].l_um_iw[205] ;
 wire \top_I.branch[11].l_um_iw[206] ;
 wire \top_I.branch[11].l_um_iw[207] ;
 wire \top_I.branch[11].l_um_iw[208] ;
 wire \top_I.branch[11].l_um_iw[209] ;
 wire \top_I.branch[11].l_um_iw[20] ;
 wire \top_I.branch[11].l_um_iw[210] ;
 wire \top_I.branch[11].l_um_iw[211] ;
 wire \top_I.branch[11].l_um_iw[212] ;
 wire \top_I.branch[11].l_um_iw[213] ;
 wire \top_I.branch[11].l_um_iw[214] ;
 wire \top_I.branch[11].l_um_iw[215] ;
 wire \top_I.branch[11].l_um_iw[216] ;
 wire \top_I.branch[11].l_um_iw[217] ;
 wire \top_I.branch[11].l_um_iw[218] ;
 wire \top_I.branch[11].l_um_iw[219] ;
 wire \top_I.branch[11].l_um_iw[21] ;
 wire \top_I.branch[11].l_um_iw[220] ;
 wire \top_I.branch[11].l_um_iw[221] ;
 wire \top_I.branch[11].l_um_iw[222] ;
 wire \top_I.branch[11].l_um_iw[223] ;
 wire \top_I.branch[11].l_um_iw[224] ;
 wire \top_I.branch[11].l_um_iw[225] ;
 wire \top_I.branch[11].l_um_iw[226] ;
 wire \top_I.branch[11].l_um_iw[227] ;
 wire \top_I.branch[11].l_um_iw[228] ;
 wire \top_I.branch[11].l_um_iw[229] ;
 wire \top_I.branch[11].l_um_iw[22] ;
 wire \top_I.branch[11].l_um_iw[230] ;
 wire \top_I.branch[11].l_um_iw[231] ;
 wire \top_I.branch[11].l_um_iw[232] ;
 wire \top_I.branch[11].l_um_iw[233] ;
 wire \top_I.branch[11].l_um_iw[234] ;
 wire \top_I.branch[11].l_um_iw[235] ;
 wire \top_I.branch[11].l_um_iw[236] ;
 wire \top_I.branch[11].l_um_iw[237] ;
 wire \top_I.branch[11].l_um_iw[238] ;
 wire \top_I.branch[11].l_um_iw[239] ;
 wire \top_I.branch[11].l_um_iw[23] ;
 wire \top_I.branch[11].l_um_iw[240] ;
 wire \top_I.branch[11].l_um_iw[241] ;
 wire \top_I.branch[11].l_um_iw[242] ;
 wire \top_I.branch[11].l_um_iw[243] ;
 wire \top_I.branch[11].l_um_iw[244] ;
 wire \top_I.branch[11].l_um_iw[245] ;
 wire \top_I.branch[11].l_um_iw[246] ;
 wire \top_I.branch[11].l_um_iw[247] ;
 wire \top_I.branch[11].l_um_iw[248] ;
 wire \top_I.branch[11].l_um_iw[249] ;
 wire \top_I.branch[11].l_um_iw[24] ;
 wire \top_I.branch[11].l_um_iw[250] ;
 wire \top_I.branch[11].l_um_iw[251] ;
 wire \top_I.branch[11].l_um_iw[252] ;
 wire \top_I.branch[11].l_um_iw[253] ;
 wire \top_I.branch[11].l_um_iw[254] ;
 wire \top_I.branch[11].l_um_iw[255] ;
 wire \top_I.branch[11].l_um_iw[256] ;
 wire \top_I.branch[11].l_um_iw[257] ;
 wire \top_I.branch[11].l_um_iw[258] ;
 wire \top_I.branch[11].l_um_iw[259] ;
 wire \top_I.branch[11].l_um_iw[25] ;
 wire \top_I.branch[11].l_um_iw[260] ;
 wire \top_I.branch[11].l_um_iw[261] ;
 wire \top_I.branch[11].l_um_iw[262] ;
 wire \top_I.branch[11].l_um_iw[263] ;
 wire \top_I.branch[11].l_um_iw[264] ;
 wire \top_I.branch[11].l_um_iw[265] ;
 wire \top_I.branch[11].l_um_iw[266] ;
 wire \top_I.branch[11].l_um_iw[267] ;
 wire \top_I.branch[11].l_um_iw[268] ;
 wire \top_I.branch[11].l_um_iw[269] ;
 wire \top_I.branch[11].l_um_iw[26] ;
 wire \top_I.branch[11].l_um_iw[270] ;
 wire \top_I.branch[11].l_um_iw[271] ;
 wire \top_I.branch[11].l_um_iw[272] ;
 wire \top_I.branch[11].l_um_iw[273] ;
 wire \top_I.branch[11].l_um_iw[274] ;
 wire \top_I.branch[11].l_um_iw[275] ;
 wire \top_I.branch[11].l_um_iw[276] ;
 wire \top_I.branch[11].l_um_iw[277] ;
 wire \top_I.branch[11].l_um_iw[278] ;
 wire \top_I.branch[11].l_um_iw[279] ;
 wire \top_I.branch[11].l_um_iw[27] ;
 wire \top_I.branch[11].l_um_iw[280] ;
 wire \top_I.branch[11].l_um_iw[281] ;
 wire \top_I.branch[11].l_um_iw[282] ;
 wire \top_I.branch[11].l_um_iw[283] ;
 wire \top_I.branch[11].l_um_iw[284] ;
 wire \top_I.branch[11].l_um_iw[285] ;
 wire \top_I.branch[11].l_um_iw[286] ;
 wire \top_I.branch[11].l_um_iw[287] ;
 wire \top_I.branch[11].l_um_iw[28] ;
 wire \top_I.branch[11].l_um_iw[29] ;
 wire \top_I.branch[11].l_um_iw[2] ;
 wire \top_I.branch[11].l_um_iw[30] ;
 wire \top_I.branch[11].l_um_iw[31] ;
 wire \top_I.branch[11].l_um_iw[32] ;
 wire \top_I.branch[11].l_um_iw[33] ;
 wire \top_I.branch[11].l_um_iw[34] ;
 wire \top_I.branch[11].l_um_iw[35] ;
 wire \top_I.branch[11].l_um_iw[36] ;
 wire \top_I.branch[11].l_um_iw[37] ;
 wire \top_I.branch[11].l_um_iw[38] ;
 wire \top_I.branch[11].l_um_iw[39] ;
 wire \top_I.branch[11].l_um_iw[3] ;
 wire \top_I.branch[11].l_um_iw[40] ;
 wire \top_I.branch[11].l_um_iw[41] ;
 wire \top_I.branch[11].l_um_iw[42] ;
 wire \top_I.branch[11].l_um_iw[43] ;
 wire \top_I.branch[11].l_um_iw[44] ;
 wire \top_I.branch[11].l_um_iw[45] ;
 wire \top_I.branch[11].l_um_iw[46] ;
 wire \top_I.branch[11].l_um_iw[47] ;
 wire \top_I.branch[11].l_um_iw[48] ;
 wire \top_I.branch[11].l_um_iw[49] ;
 wire \top_I.branch[11].l_um_iw[4] ;
 wire \top_I.branch[11].l_um_iw[50] ;
 wire \top_I.branch[11].l_um_iw[51] ;
 wire \top_I.branch[11].l_um_iw[52] ;
 wire \top_I.branch[11].l_um_iw[53] ;
 wire \top_I.branch[11].l_um_iw[54] ;
 wire \top_I.branch[11].l_um_iw[55] ;
 wire \top_I.branch[11].l_um_iw[56] ;
 wire \top_I.branch[11].l_um_iw[57] ;
 wire \top_I.branch[11].l_um_iw[58] ;
 wire \top_I.branch[11].l_um_iw[59] ;
 wire \top_I.branch[11].l_um_iw[5] ;
 wire \top_I.branch[11].l_um_iw[60] ;
 wire \top_I.branch[11].l_um_iw[61] ;
 wire \top_I.branch[11].l_um_iw[62] ;
 wire \top_I.branch[11].l_um_iw[63] ;
 wire \top_I.branch[11].l_um_iw[64] ;
 wire \top_I.branch[11].l_um_iw[65] ;
 wire \top_I.branch[11].l_um_iw[66] ;
 wire \top_I.branch[11].l_um_iw[67] ;
 wire \top_I.branch[11].l_um_iw[68] ;
 wire \top_I.branch[11].l_um_iw[69] ;
 wire \top_I.branch[11].l_um_iw[6] ;
 wire \top_I.branch[11].l_um_iw[70] ;
 wire \top_I.branch[11].l_um_iw[71] ;
 wire \top_I.branch[11].l_um_iw[72] ;
 wire \top_I.branch[11].l_um_iw[73] ;
 wire \top_I.branch[11].l_um_iw[74] ;
 wire \top_I.branch[11].l_um_iw[75] ;
 wire \top_I.branch[11].l_um_iw[76] ;
 wire \top_I.branch[11].l_um_iw[77] ;
 wire \top_I.branch[11].l_um_iw[78] ;
 wire \top_I.branch[11].l_um_iw[79] ;
 wire \top_I.branch[11].l_um_iw[7] ;
 wire \top_I.branch[11].l_um_iw[80] ;
 wire \top_I.branch[11].l_um_iw[81] ;
 wire \top_I.branch[11].l_um_iw[82] ;
 wire \top_I.branch[11].l_um_iw[83] ;
 wire \top_I.branch[11].l_um_iw[84] ;
 wire \top_I.branch[11].l_um_iw[85] ;
 wire \top_I.branch[11].l_um_iw[86] ;
 wire \top_I.branch[11].l_um_iw[87] ;
 wire \top_I.branch[11].l_um_iw[88] ;
 wire \top_I.branch[11].l_um_iw[89] ;
 wire \top_I.branch[11].l_um_iw[8] ;
 wire \top_I.branch[11].l_um_iw[90] ;
 wire \top_I.branch[11].l_um_iw[91] ;
 wire \top_I.branch[11].l_um_iw[92] ;
 wire \top_I.branch[11].l_um_iw[93] ;
 wire \top_I.branch[11].l_um_iw[94] ;
 wire \top_I.branch[11].l_um_iw[95] ;
 wire \top_I.branch[11].l_um_iw[96] ;
 wire \top_I.branch[11].l_um_iw[97] ;
 wire \top_I.branch[11].l_um_iw[98] ;
 wire \top_I.branch[11].l_um_iw[99] ;
 wire \top_I.branch[11].l_um_iw[9] ;
 wire \top_I.branch[11].l_um_k_zero[0] ;
 wire \top_I.branch[11].l_um_k_zero[10] ;
 wire \top_I.branch[11].l_um_k_zero[11] ;
 wire \top_I.branch[11].l_um_k_zero[12] ;
 wire \top_I.branch[11].l_um_k_zero[13] ;
 wire \top_I.branch[11].l_um_k_zero[14] ;
 wire \top_I.branch[11].l_um_k_zero[15] ;
 wire \top_I.branch[11].l_um_k_zero[1] ;
 wire \top_I.branch[11].l_um_k_zero[2] ;
 wire \top_I.branch[11].l_um_k_zero[3] ;
 wire \top_I.branch[11].l_um_k_zero[4] ;
 wire \top_I.branch[11].l_um_k_zero[5] ;
 wire \top_I.branch[11].l_um_k_zero[6] ;
 wire \top_I.branch[11].l_um_k_zero[7] ;
 wire \top_I.branch[11].l_um_k_zero[8] ;
 wire \top_I.branch[11].l_um_k_zero[9] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[12].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[12].l_k_one ;
 wire \top_I.branch[12].l_k_zero ;
 wire \top_I.branch[12].l_um_ena[0] ;
 wire \top_I.branch[12].l_um_ena[10] ;
 wire \top_I.branch[12].l_um_ena[11] ;
 wire \top_I.branch[12].l_um_ena[12] ;
 wire \top_I.branch[12].l_um_ena[13] ;
 wire \top_I.branch[12].l_um_ena[14] ;
 wire \top_I.branch[12].l_um_ena[15] ;
 wire \top_I.branch[12].l_um_ena[1] ;
 wire \top_I.branch[12].l_um_ena[2] ;
 wire \top_I.branch[12].l_um_ena[3] ;
 wire \top_I.branch[12].l_um_ena[4] ;
 wire \top_I.branch[12].l_um_ena[5] ;
 wire \top_I.branch[12].l_um_ena[6] ;
 wire \top_I.branch[12].l_um_ena[7] ;
 wire \top_I.branch[12].l_um_ena[8] ;
 wire \top_I.branch[12].l_um_ena[9] ;
 wire \top_I.branch[12].l_um_iw[0] ;
 wire \top_I.branch[12].l_um_iw[100] ;
 wire \top_I.branch[12].l_um_iw[101] ;
 wire \top_I.branch[12].l_um_iw[102] ;
 wire \top_I.branch[12].l_um_iw[103] ;
 wire \top_I.branch[12].l_um_iw[104] ;
 wire \top_I.branch[12].l_um_iw[105] ;
 wire \top_I.branch[12].l_um_iw[106] ;
 wire \top_I.branch[12].l_um_iw[107] ;
 wire \top_I.branch[12].l_um_iw[108] ;
 wire \top_I.branch[12].l_um_iw[109] ;
 wire \top_I.branch[12].l_um_iw[10] ;
 wire \top_I.branch[12].l_um_iw[110] ;
 wire \top_I.branch[12].l_um_iw[111] ;
 wire \top_I.branch[12].l_um_iw[112] ;
 wire \top_I.branch[12].l_um_iw[113] ;
 wire \top_I.branch[12].l_um_iw[114] ;
 wire \top_I.branch[12].l_um_iw[115] ;
 wire \top_I.branch[12].l_um_iw[116] ;
 wire \top_I.branch[12].l_um_iw[117] ;
 wire \top_I.branch[12].l_um_iw[118] ;
 wire \top_I.branch[12].l_um_iw[119] ;
 wire \top_I.branch[12].l_um_iw[11] ;
 wire \top_I.branch[12].l_um_iw[120] ;
 wire \top_I.branch[12].l_um_iw[121] ;
 wire \top_I.branch[12].l_um_iw[122] ;
 wire \top_I.branch[12].l_um_iw[123] ;
 wire \top_I.branch[12].l_um_iw[124] ;
 wire \top_I.branch[12].l_um_iw[125] ;
 wire \top_I.branch[12].l_um_iw[126] ;
 wire \top_I.branch[12].l_um_iw[127] ;
 wire \top_I.branch[12].l_um_iw[128] ;
 wire \top_I.branch[12].l_um_iw[129] ;
 wire \top_I.branch[12].l_um_iw[12] ;
 wire \top_I.branch[12].l_um_iw[130] ;
 wire \top_I.branch[12].l_um_iw[131] ;
 wire \top_I.branch[12].l_um_iw[132] ;
 wire \top_I.branch[12].l_um_iw[133] ;
 wire \top_I.branch[12].l_um_iw[134] ;
 wire \top_I.branch[12].l_um_iw[135] ;
 wire \top_I.branch[12].l_um_iw[136] ;
 wire \top_I.branch[12].l_um_iw[137] ;
 wire \top_I.branch[12].l_um_iw[138] ;
 wire \top_I.branch[12].l_um_iw[139] ;
 wire \top_I.branch[12].l_um_iw[13] ;
 wire \top_I.branch[12].l_um_iw[140] ;
 wire \top_I.branch[12].l_um_iw[141] ;
 wire \top_I.branch[12].l_um_iw[142] ;
 wire \top_I.branch[12].l_um_iw[143] ;
 wire \top_I.branch[12].l_um_iw[144] ;
 wire \top_I.branch[12].l_um_iw[145] ;
 wire \top_I.branch[12].l_um_iw[146] ;
 wire \top_I.branch[12].l_um_iw[147] ;
 wire \top_I.branch[12].l_um_iw[148] ;
 wire \top_I.branch[12].l_um_iw[149] ;
 wire \top_I.branch[12].l_um_iw[14] ;
 wire \top_I.branch[12].l_um_iw[150] ;
 wire \top_I.branch[12].l_um_iw[151] ;
 wire \top_I.branch[12].l_um_iw[152] ;
 wire \top_I.branch[12].l_um_iw[153] ;
 wire \top_I.branch[12].l_um_iw[154] ;
 wire \top_I.branch[12].l_um_iw[155] ;
 wire \top_I.branch[12].l_um_iw[156] ;
 wire \top_I.branch[12].l_um_iw[157] ;
 wire \top_I.branch[12].l_um_iw[158] ;
 wire \top_I.branch[12].l_um_iw[159] ;
 wire \top_I.branch[12].l_um_iw[15] ;
 wire \top_I.branch[12].l_um_iw[160] ;
 wire \top_I.branch[12].l_um_iw[161] ;
 wire \top_I.branch[12].l_um_iw[162] ;
 wire \top_I.branch[12].l_um_iw[163] ;
 wire \top_I.branch[12].l_um_iw[164] ;
 wire \top_I.branch[12].l_um_iw[165] ;
 wire \top_I.branch[12].l_um_iw[166] ;
 wire \top_I.branch[12].l_um_iw[167] ;
 wire \top_I.branch[12].l_um_iw[168] ;
 wire \top_I.branch[12].l_um_iw[169] ;
 wire \top_I.branch[12].l_um_iw[16] ;
 wire \top_I.branch[12].l_um_iw[170] ;
 wire \top_I.branch[12].l_um_iw[171] ;
 wire \top_I.branch[12].l_um_iw[172] ;
 wire \top_I.branch[12].l_um_iw[173] ;
 wire \top_I.branch[12].l_um_iw[174] ;
 wire \top_I.branch[12].l_um_iw[175] ;
 wire \top_I.branch[12].l_um_iw[176] ;
 wire \top_I.branch[12].l_um_iw[177] ;
 wire \top_I.branch[12].l_um_iw[178] ;
 wire \top_I.branch[12].l_um_iw[179] ;
 wire \top_I.branch[12].l_um_iw[17] ;
 wire \top_I.branch[12].l_um_iw[180] ;
 wire \top_I.branch[12].l_um_iw[181] ;
 wire \top_I.branch[12].l_um_iw[182] ;
 wire \top_I.branch[12].l_um_iw[183] ;
 wire \top_I.branch[12].l_um_iw[184] ;
 wire \top_I.branch[12].l_um_iw[185] ;
 wire \top_I.branch[12].l_um_iw[186] ;
 wire \top_I.branch[12].l_um_iw[187] ;
 wire \top_I.branch[12].l_um_iw[188] ;
 wire \top_I.branch[12].l_um_iw[189] ;
 wire \top_I.branch[12].l_um_iw[18] ;
 wire \top_I.branch[12].l_um_iw[190] ;
 wire \top_I.branch[12].l_um_iw[191] ;
 wire \top_I.branch[12].l_um_iw[192] ;
 wire \top_I.branch[12].l_um_iw[193] ;
 wire \top_I.branch[12].l_um_iw[194] ;
 wire \top_I.branch[12].l_um_iw[195] ;
 wire \top_I.branch[12].l_um_iw[196] ;
 wire \top_I.branch[12].l_um_iw[197] ;
 wire \top_I.branch[12].l_um_iw[198] ;
 wire \top_I.branch[12].l_um_iw[199] ;
 wire \top_I.branch[12].l_um_iw[19] ;
 wire \top_I.branch[12].l_um_iw[1] ;
 wire \top_I.branch[12].l_um_iw[200] ;
 wire \top_I.branch[12].l_um_iw[201] ;
 wire \top_I.branch[12].l_um_iw[202] ;
 wire \top_I.branch[12].l_um_iw[203] ;
 wire \top_I.branch[12].l_um_iw[204] ;
 wire \top_I.branch[12].l_um_iw[205] ;
 wire \top_I.branch[12].l_um_iw[206] ;
 wire \top_I.branch[12].l_um_iw[207] ;
 wire \top_I.branch[12].l_um_iw[208] ;
 wire \top_I.branch[12].l_um_iw[209] ;
 wire \top_I.branch[12].l_um_iw[20] ;
 wire \top_I.branch[12].l_um_iw[210] ;
 wire \top_I.branch[12].l_um_iw[211] ;
 wire \top_I.branch[12].l_um_iw[212] ;
 wire \top_I.branch[12].l_um_iw[213] ;
 wire \top_I.branch[12].l_um_iw[214] ;
 wire \top_I.branch[12].l_um_iw[215] ;
 wire \top_I.branch[12].l_um_iw[216] ;
 wire \top_I.branch[12].l_um_iw[217] ;
 wire \top_I.branch[12].l_um_iw[218] ;
 wire \top_I.branch[12].l_um_iw[219] ;
 wire \top_I.branch[12].l_um_iw[21] ;
 wire \top_I.branch[12].l_um_iw[220] ;
 wire \top_I.branch[12].l_um_iw[221] ;
 wire \top_I.branch[12].l_um_iw[222] ;
 wire \top_I.branch[12].l_um_iw[223] ;
 wire \top_I.branch[12].l_um_iw[224] ;
 wire \top_I.branch[12].l_um_iw[225] ;
 wire \top_I.branch[12].l_um_iw[226] ;
 wire \top_I.branch[12].l_um_iw[227] ;
 wire \top_I.branch[12].l_um_iw[228] ;
 wire \top_I.branch[12].l_um_iw[229] ;
 wire \top_I.branch[12].l_um_iw[22] ;
 wire \top_I.branch[12].l_um_iw[230] ;
 wire \top_I.branch[12].l_um_iw[231] ;
 wire \top_I.branch[12].l_um_iw[232] ;
 wire \top_I.branch[12].l_um_iw[233] ;
 wire \top_I.branch[12].l_um_iw[234] ;
 wire \top_I.branch[12].l_um_iw[235] ;
 wire \top_I.branch[12].l_um_iw[236] ;
 wire \top_I.branch[12].l_um_iw[237] ;
 wire \top_I.branch[12].l_um_iw[238] ;
 wire \top_I.branch[12].l_um_iw[239] ;
 wire \top_I.branch[12].l_um_iw[23] ;
 wire \top_I.branch[12].l_um_iw[240] ;
 wire \top_I.branch[12].l_um_iw[241] ;
 wire \top_I.branch[12].l_um_iw[242] ;
 wire \top_I.branch[12].l_um_iw[243] ;
 wire \top_I.branch[12].l_um_iw[244] ;
 wire \top_I.branch[12].l_um_iw[245] ;
 wire \top_I.branch[12].l_um_iw[246] ;
 wire \top_I.branch[12].l_um_iw[247] ;
 wire \top_I.branch[12].l_um_iw[248] ;
 wire \top_I.branch[12].l_um_iw[249] ;
 wire \top_I.branch[12].l_um_iw[24] ;
 wire \top_I.branch[12].l_um_iw[250] ;
 wire \top_I.branch[12].l_um_iw[251] ;
 wire \top_I.branch[12].l_um_iw[252] ;
 wire \top_I.branch[12].l_um_iw[253] ;
 wire \top_I.branch[12].l_um_iw[254] ;
 wire \top_I.branch[12].l_um_iw[255] ;
 wire \top_I.branch[12].l_um_iw[256] ;
 wire \top_I.branch[12].l_um_iw[257] ;
 wire \top_I.branch[12].l_um_iw[258] ;
 wire \top_I.branch[12].l_um_iw[259] ;
 wire \top_I.branch[12].l_um_iw[25] ;
 wire \top_I.branch[12].l_um_iw[260] ;
 wire \top_I.branch[12].l_um_iw[261] ;
 wire \top_I.branch[12].l_um_iw[262] ;
 wire \top_I.branch[12].l_um_iw[263] ;
 wire \top_I.branch[12].l_um_iw[264] ;
 wire \top_I.branch[12].l_um_iw[265] ;
 wire \top_I.branch[12].l_um_iw[266] ;
 wire \top_I.branch[12].l_um_iw[267] ;
 wire \top_I.branch[12].l_um_iw[268] ;
 wire \top_I.branch[12].l_um_iw[269] ;
 wire \top_I.branch[12].l_um_iw[26] ;
 wire \top_I.branch[12].l_um_iw[270] ;
 wire \top_I.branch[12].l_um_iw[271] ;
 wire \top_I.branch[12].l_um_iw[272] ;
 wire \top_I.branch[12].l_um_iw[273] ;
 wire \top_I.branch[12].l_um_iw[274] ;
 wire \top_I.branch[12].l_um_iw[275] ;
 wire \top_I.branch[12].l_um_iw[276] ;
 wire \top_I.branch[12].l_um_iw[277] ;
 wire \top_I.branch[12].l_um_iw[278] ;
 wire \top_I.branch[12].l_um_iw[279] ;
 wire \top_I.branch[12].l_um_iw[27] ;
 wire \top_I.branch[12].l_um_iw[280] ;
 wire \top_I.branch[12].l_um_iw[281] ;
 wire \top_I.branch[12].l_um_iw[282] ;
 wire \top_I.branch[12].l_um_iw[283] ;
 wire \top_I.branch[12].l_um_iw[284] ;
 wire \top_I.branch[12].l_um_iw[285] ;
 wire \top_I.branch[12].l_um_iw[286] ;
 wire \top_I.branch[12].l_um_iw[287] ;
 wire \top_I.branch[12].l_um_iw[28] ;
 wire \top_I.branch[12].l_um_iw[29] ;
 wire \top_I.branch[12].l_um_iw[2] ;
 wire \top_I.branch[12].l_um_iw[30] ;
 wire \top_I.branch[12].l_um_iw[31] ;
 wire \top_I.branch[12].l_um_iw[32] ;
 wire \top_I.branch[12].l_um_iw[33] ;
 wire \top_I.branch[12].l_um_iw[34] ;
 wire \top_I.branch[12].l_um_iw[35] ;
 wire \top_I.branch[12].l_um_iw[36] ;
 wire \top_I.branch[12].l_um_iw[37] ;
 wire \top_I.branch[12].l_um_iw[38] ;
 wire \top_I.branch[12].l_um_iw[39] ;
 wire \top_I.branch[12].l_um_iw[3] ;
 wire \top_I.branch[12].l_um_iw[40] ;
 wire \top_I.branch[12].l_um_iw[41] ;
 wire \top_I.branch[12].l_um_iw[42] ;
 wire \top_I.branch[12].l_um_iw[43] ;
 wire \top_I.branch[12].l_um_iw[44] ;
 wire \top_I.branch[12].l_um_iw[45] ;
 wire \top_I.branch[12].l_um_iw[46] ;
 wire \top_I.branch[12].l_um_iw[47] ;
 wire \top_I.branch[12].l_um_iw[48] ;
 wire \top_I.branch[12].l_um_iw[49] ;
 wire \top_I.branch[12].l_um_iw[4] ;
 wire \top_I.branch[12].l_um_iw[50] ;
 wire \top_I.branch[12].l_um_iw[51] ;
 wire \top_I.branch[12].l_um_iw[52] ;
 wire \top_I.branch[12].l_um_iw[53] ;
 wire \top_I.branch[12].l_um_iw[54] ;
 wire \top_I.branch[12].l_um_iw[55] ;
 wire \top_I.branch[12].l_um_iw[56] ;
 wire \top_I.branch[12].l_um_iw[57] ;
 wire \top_I.branch[12].l_um_iw[58] ;
 wire \top_I.branch[12].l_um_iw[59] ;
 wire \top_I.branch[12].l_um_iw[5] ;
 wire \top_I.branch[12].l_um_iw[60] ;
 wire \top_I.branch[12].l_um_iw[61] ;
 wire \top_I.branch[12].l_um_iw[62] ;
 wire \top_I.branch[12].l_um_iw[63] ;
 wire \top_I.branch[12].l_um_iw[64] ;
 wire \top_I.branch[12].l_um_iw[65] ;
 wire \top_I.branch[12].l_um_iw[66] ;
 wire \top_I.branch[12].l_um_iw[67] ;
 wire \top_I.branch[12].l_um_iw[68] ;
 wire \top_I.branch[12].l_um_iw[69] ;
 wire \top_I.branch[12].l_um_iw[6] ;
 wire \top_I.branch[12].l_um_iw[70] ;
 wire \top_I.branch[12].l_um_iw[71] ;
 wire \top_I.branch[12].l_um_iw[72] ;
 wire \top_I.branch[12].l_um_iw[73] ;
 wire \top_I.branch[12].l_um_iw[74] ;
 wire \top_I.branch[12].l_um_iw[75] ;
 wire \top_I.branch[12].l_um_iw[76] ;
 wire \top_I.branch[12].l_um_iw[77] ;
 wire \top_I.branch[12].l_um_iw[78] ;
 wire \top_I.branch[12].l_um_iw[79] ;
 wire \top_I.branch[12].l_um_iw[7] ;
 wire \top_I.branch[12].l_um_iw[80] ;
 wire \top_I.branch[12].l_um_iw[81] ;
 wire \top_I.branch[12].l_um_iw[82] ;
 wire \top_I.branch[12].l_um_iw[83] ;
 wire \top_I.branch[12].l_um_iw[84] ;
 wire \top_I.branch[12].l_um_iw[85] ;
 wire \top_I.branch[12].l_um_iw[86] ;
 wire \top_I.branch[12].l_um_iw[87] ;
 wire \top_I.branch[12].l_um_iw[88] ;
 wire \top_I.branch[12].l_um_iw[89] ;
 wire \top_I.branch[12].l_um_iw[8] ;
 wire \top_I.branch[12].l_um_iw[90] ;
 wire \top_I.branch[12].l_um_iw[91] ;
 wire \top_I.branch[12].l_um_iw[92] ;
 wire \top_I.branch[12].l_um_iw[93] ;
 wire \top_I.branch[12].l_um_iw[94] ;
 wire \top_I.branch[12].l_um_iw[95] ;
 wire \top_I.branch[12].l_um_iw[96] ;
 wire \top_I.branch[12].l_um_iw[97] ;
 wire \top_I.branch[12].l_um_iw[98] ;
 wire \top_I.branch[12].l_um_iw[99] ;
 wire \top_I.branch[12].l_um_iw[9] ;
 wire \top_I.branch[12].l_um_k_zero[0] ;
 wire \top_I.branch[12].l_um_k_zero[10] ;
 wire \top_I.branch[12].l_um_k_zero[11] ;
 wire \top_I.branch[12].l_um_k_zero[12] ;
 wire \top_I.branch[12].l_um_k_zero[13] ;
 wire \top_I.branch[12].l_um_k_zero[14] ;
 wire \top_I.branch[12].l_um_k_zero[15] ;
 wire \top_I.branch[12].l_um_k_zero[1] ;
 wire \top_I.branch[12].l_um_k_zero[2] ;
 wire \top_I.branch[12].l_um_k_zero[3] ;
 wire \top_I.branch[12].l_um_k_zero[4] ;
 wire \top_I.branch[12].l_um_k_zero[5] ;
 wire \top_I.branch[12].l_um_k_zero[6] ;
 wire \top_I.branch[12].l_um_k_zero[7] ;
 wire \top_I.branch[12].l_um_k_zero[8] ;
 wire \top_I.branch[12].l_um_k_zero[9] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[13].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[13].l_k_one ;
 wire \top_I.branch[13].l_k_zero ;
 wire \top_I.branch[13].l_um_ena[0] ;
 wire \top_I.branch[13].l_um_ena[10] ;
 wire \top_I.branch[13].l_um_ena[11] ;
 wire \top_I.branch[13].l_um_ena[12] ;
 wire \top_I.branch[13].l_um_ena[13] ;
 wire \top_I.branch[13].l_um_ena[14] ;
 wire \top_I.branch[13].l_um_ena[15] ;
 wire \top_I.branch[13].l_um_ena[1] ;
 wire \top_I.branch[13].l_um_ena[2] ;
 wire \top_I.branch[13].l_um_ena[3] ;
 wire \top_I.branch[13].l_um_ena[4] ;
 wire \top_I.branch[13].l_um_ena[5] ;
 wire \top_I.branch[13].l_um_ena[6] ;
 wire \top_I.branch[13].l_um_ena[7] ;
 wire \top_I.branch[13].l_um_ena[8] ;
 wire \top_I.branch[13].l_um_ena[9] ;
 wire \top_I.branch[13].l_um_iw[0] ;
 wire \top_I.branch[13].l_um_iw[100] ;
 wire \top_I.branch[13].l_um_iw[101] ;
 wire \top_I.branch[13].l_um_iw[102] ;
 wire \top_I.branch[13].l_um_iw[103] ;
 wire \top_I.branch[13].l_um_iw[104] ;
 wire \top_I.branch[13].l_um_iw[105] ;
 wire \top_I.branch[13].l_um_iw[106] ;
 wire \top_I.branch[13].l_um_iw[107] ;
 wire \top_I.branch[13].l_um_iw[108] ;
 wire \top_I.branch[13].l_um_iw[109] ;
 wire \top_I.branch[13].l_um_iw[10] ;
 wire \top_I.branch[13].l_um_iw[110] ;
 wire \top_I.branch[13].l_um_iw[111] ;
 wire \top_I.branch[13].l_um_iw[112] ;
 wire \top_I.branch[13].l_um_iw[113] ;
 wire \top_I.branch[13].l_um_iw[114] ;
 wire \top_I.branch[13].l_um_iw[115] ;
 wire \top_I.branch[13].l_um_iw[116] ;
 wire \top_I.branch[13].l_um_iw[117] ;
 wire \top_I.branch[13].l_um_iw[118] ;
 wire \top_I.branch[13].l_um_iw[119] ;
 wire \top_I.branch[13].l_um_iw[11] ;
 wire \top_I.branch[13].l_um_iw[120] ;
 wire \top_I.branch[13].l_um_iw[121] ;
 wire \top_I.branch[13].l_um_iw[122] ;
 wire \top_I.branch[13].l_um_iw[123] ;
 wire \top_I.branch[13].l_um_iw[124] ;
 wire \top_I.branch[13].l_um_iw[125] ;
 wire \top_I.branch[13].l_um_iw[126] ;
 wire \top_I.branch[13].l_um_iw[127] ;
 wire \top_I.branch[13].l_um_iw[128] ;
 wire \top_I.branch[13].l_um_iw[129] ;
 wire \top_I.branch[13].l_um_iw[12] ;
 wire \top_I.branch[13].l_um_iw[130] ;
 wire \top_I.branch[13].l_um_iw[131] ;
 wire \top_I.branch[13].l_um_iw[132] ;
 wire \top_I.branch[13].l_um_iw[133] ;
 wire \top_I.branch[13].l_um_iw[134] ;
 wire \top_I.branch[13].l_um_iw[135] ;
 wire \top_I.branch[13].l_um_iw[136] ;
 wire \top_I.branch[13].l_um_iw[137] ;
 wire \top_I.branch[13].l_um_iw[138] ;
 wire \top_I.branch[13].l_um_iw[139] ;
 wire \top_I.branch[13].l_um_iw[13] ;
 wire \top_I.branch[13].l_um_iw[140] ;
 wire \top_I.branch[13].l_um_iw[141] ;
 wire \top_I.branch[13].l_um_iw[142] ;
 wire \top_I.branch[13].l_um_iw[143] ;
 wire \top_I.branch[13].l_um_iw[144] ;
 wire \top_I.branch[13].l_um_iw[145] ;
 wire \top_I.branch[13].l_um_iw[146] ;
 wire \top_I.branch[13].l_um_iw[147] ;
 wire \top_I.branch[13].l_um_iw[148] ;
 wire \top_I.branch[13].l_um_iw[149] ;
 wire \top_I.branch[13].l_um_iw[14] ;
 wire \top_I.branch[13].l_um_iw[150] ;
 wire \top_I.branch[13].l_um_iw[151] ;
 wire \top_I.branch[13].l_um_iw[152] ;
 wire \top_I.branch[13].l_um_iw[153] ;
 wire \top_I.branch[13].l_um_iw[154] ;
 wire \top_I.branch[13].l_um_iw[155] ;
 wire \top_I.branch[13].l_um_iw[156] ;
 wire \top_I.branch[13].l_um_iw[157] ;
 wire \top_I.branch[13].l_um_iw[158] ;
 wire \top_I.branch[13].l_um_iw[159] ;
 wire \top_I.branch[13].l_um_iw[15] ;
 wire \top_I.branch[13].l_um_iw[160] ;
 wire \top_I.branch[13].l_um_iw[161] ;
 wire \top_I.branch[13].l_um_iw[162] ;
 wire \top_I.branch[13].l_um_iw[163] ;
 wire \top_I.branch[13].l_um_iw[164] ;
 wire \top_I.branch[13].l_um_iw[165] ;
 wire \top_I.branch[13].l_um_iw[166] ;
 wire \top_I.branch[13].l_um_iw[167] ;
 wire \top_I.branch[13].l_um_iw[168] ;
 wire \top_I.branch[13].l_um_iw[169] ;
 wire \top_I.branch[13].l_um_iw[16] ;
 wire \top_I.branch[13].l_um_iw[170] ;
 wire \top_I.branch[13].l_um_iw[171] ;
 wire \top_I.branch[13].l_um_iw[172] ;
 wire \top_I.branch[13].l_um_iw[173] ;
 wire \top_I.branch[13].l_um_iw[174] ;
 wire \top_I.branch[13].l_um_iw[175] ;
 wire \top_I.branch[13].l_um_iw[176] ;
 wire \top_I.branch[13].l_um_iw[177] ;
 wire \top_I.branch[13].l_um_iw[178] ;
 wire \top_I.branch[13].l_um_iw[179] ;
 wire \top_I.branch[13].l_um_iw[17] ;
 wire \top_I.branch[13].l_um_iw[180] ;
 wire \top_I.branch[13].l_um_iw[181] ;
 wire \top_I.branch[13].l_um_iw[182] ;
 wire \top_I.branch[13].l_um_iw[183] ;
 wire \top_I.branch[13].l_um_iw[184] ;
 wire \top_I.branch[13].l_um_iw[185] ;
 wire \top_I.branch[13].l_um_iw[186] ;
 wire \top_I.branch[13].l_um_iw[187] ;
 wire \top_I.branch[13].l_um_iw[188] ;
 wire \top_I.branch[13].l_um_iw[189] ;
 wire \top_I.branch[13].l_um_iw[18] ;
 wire \top_I.branch[13].l_um_iw[190] ;
 wire \top_I.branch[13].l_um_iw[191] ;
 wire \top_I.branch[13].l_um_iw[192] ;
 wire \top_I.branch[13].l_um_iw[193] ;
 wire \top_I.branch[13].l_um_iw[194] ;
 wire \top_I.branch[13].l_um_iw[195] ;
 wire \top_I.branch[13].l_um_iw[196] ;
 wire \top_I.branch[13].l_um_iw[197] ;
 wire \top_I.branch[13].l_um_iw[198] ;
 wire \top_I.branch[13].l_um_iw[199] ;
 wire \top_I.branch[13].l_um_iw[19] ;
 wire \top_I.branch[13].l_um_iw[1] ;
 wire \top_I.branch[13].l_um_iw[200] ;
 wire \top_I.branch[13].l_um_iw[201] ;
 wire \top_I.branch[13].l_um_iw[202] ;
 wire \top_I.branch[13].l_um_iw[203] ;
 wire \top_I.branch[13].l_um_iw[204] ;
 wire \top_I.branch[13].l_um_iw[205] ;
 wire \top_I.branch[13].l_um_iw[206] ;
 wire \top_I.branch[13].l_um_iw[207] ;
 wire \top_I.branch[13].l_um_iw[208] ;
 wire \top_I.branch[13].l_um_iw[209] ;
 wire \top_I.branch[13].l_um_iw[20] ;
 wire \top_I.branch[13].l_um_iw[210] ;
 wire \top_I.branch[13].l_um_iw[211] ;
 wire \top_I.branch[13].l_um_iw[212] ;
 wire \top_I.branch[13].l_um_iw[213] ;
 wire \top_I.branch[13].l_um_iw[214] ;
 wire \top_I.branch[13].l_um_iw[215] ;
 wire \top_I.branch[13].l_um_iw[216] ;
 wire \top_I.branch[13].l_um_iw[217] ;
 wire \top_I.branch[13].l_um_iw[218] ;
 wire \top_I.branch[13].l_um_iw[219] ;
 wire \top_I.branch[13].l_um_iw[21] ;
 wire \top_I.branch[13].l_um_iw[220] ;
 wire \top_I.branch[13].l_um_iw[221] ;
 wire \top_I.branch[13].l_um_iw[222] ;
 wire \top_I.branch[13].l_um_iw[223] ;
 wire \top_I.branch[13].l_um_iw[224] ;
 wire \top_I.branch[13].l_um_iw[225] ;
 wire \top_I.branch[13].l_um_iw[226] ;
 wire \top_I.branch[13].l_um_iw[227] ;
 wire \top_I.branch[13].l_um_iw[228] ;
 wire \top_I.branch[13].l_um_iw[229] ;
 wire \top_I.branch[13].l_um_iw[22] ;
 wire \top_I.branch[13].l_um_iw[230] ;
 wire \top_I.branch[13].l_um_iw[231] ;
 wire \top_I.branch[13].l_um_iw[232] ;
 wire \top_I.branch[13].l_um_iw[233] ;
 wire \top_I.branch[13].l_um_iw[234] ;
 wire \top_I.branch[13].l_um_iw[235] ;
 wire \top_I.branch[13].l_um_iw[236] ;
 wire \top_I.branch[13].l_um_iw[237] ;
 wire \top_I.branch[13].l_um_iw[238] ;
 wire \top_I.branch[13].l_um_iw[239] ;
 wire \top_I.branch[13].l_um_iw[23] ;
 wire \top_I.branch[13].l_um_iw[240] ;
 wire \top_I.branch[13].l_um_iw[241] ;
 wire \top_I.branch[13].l_um_iw[242] ;
 wire \top_I.branch[13].l_um_iw[243] ;
 wire \top_I.branch[13].l_um_iw[244] ;
 wire \top_I.branch[13].l_um_iw[245] ;
 wire \top_I.branch[13].l_um_iw[246] ;
 wire \top_I.branch[13].l_um_iw[247] ;
 wire \top_I.branch[13].l_um_iw[248] ;
 wire \top_I.branch[13].l_um_iw[249] ;
 wire \top_I.branch[13].l_um_iw[24] ;
 wire \top_I.branch[13].l_um_iw[250] ;
 wire \top_I.branch[13].l_um_iw[251] ;
 wire \top_I.branch[13].l_um_iw[252] ;
 wire \top_I.branch[13].l_um_iw[253] ;
 wire \top_I.branch[13].l_um_iw[254] ;
 wire \top_I.branch[13].l_um_iw[255] ;
 wire \top_I.branch[13].l_um_iw[256] ;
 wire \top_I.branch[13].l_um_iw[257] ;
 wire \top_I.branch[13].l_um_iw[258] ;
 wire \top_I.branch[13].l_um_iw[259] ;
 wire \top_I.branch[13].l_um_iw[25] ;
 wire \top_I.branch[13].l_um_iw[260] ;
 wire \top_I.branch[13].l_um_iw[261] ;
 wire \top_I.branch[13].l_um_iw[262] ;
 wire \top_I.branch[13].l_um_iw[263] ;
 wire \top_I.branch[13].l_um_iw[264] ;
 wire \top_I.branch[13].l_um_iw[265] ;
 wire \top_I.branch[13].l_um_iw[266] ;
 wire \top_I.branch[13].l_um_iw[267] ;
 wire \top_I.branch[13].l_um_iw[268] ;
 wire \top_I.branch[13].l_um_iw[269] ;
 wire \top_I.branch[13].l_um_iw[26] ;
 wire \top_I.branch[13].l_um_iw[270] ;
 wire \top_I.branch[13].l_um_iw[271] ;
 wire \top_I.branch[13].l_um_iw[272] ;
 wire \top_I.branch[13].l_um_iw[273] ;
 wire \top_I.branch[13].l_um_iw[274] ;
 wire \top_I.branch[13].l_um_iw[275] ;
 wire \top_I.branch[13].l_um_iw[276] ;
 wire \top_I.branch[13].l_um_iw[277] ;
 wire \top_I.branch[13].l_um_iw[278] ;
 wire \top_I.branch[13].l_um_iw[279] ;
 wire \top_I.branch[13].l_um_iw[27] ;
 wire \top_I.branch[13].l_um_iw[280] ;
 wire \top_I.branch[13].l_um_iw[281] ;
 wire \top_I.branch[13].l_um_iw[282] ;
 wire \top_I.branch[13].l_um_iw[283] ;
 wire \top_I.branch[13].l_um_iw[284] ;
 wire \top_I.branch[13].l_um_iw[285] ;
 wire \top_I.branch[13].l_um_iw[286] ;
 wire \top_I.branch[13].l_um_iw[287] ;
 wire \top_I.branch[13].l_um_iw[28] ;
 wire \top_I.branch[13].l_um_iw[29] ;
 wire \top_I.branch[13].l_um_iw[2] ;
 wire \top_I.branch[13].l_um_iw[30] ;
 wire \top_I.branch[13].l_um_iw[31] ;
 wire \top_I.branch[13].l_um_iw[32] ;
 wire \top_I.branch[13].l_um_iw[33] ;
 wire \top_I.branch[13].l_um_iw[34] ;
 wire \top_I.branch[13].l_um_iw[35] ;
 wire \top_I.branch[13].l_um_iw[36] ;
 wire \top_I.branch[13].l_um_iw[37] ;
 wire \top_I.branch[13].l_um_iw[38] ;
 wire \top_I.branch[13].l_um_iw[39] ;
 wire \top_I.branch[13].l_um_iw[3] ;
 wire \top_I.branch[13].l_um_iw[40] ;
 wire \top_I.branch[13].l_um_iw[41] ;
 wire \top_I.branch[13].l_um_iw[42] ;
 wire \top_I.branch[13].l_um_iw[43] ;
 wire \top_I.branch[13].l_um_iw[44] ;
 wire \top_I.branch[13].l_um_iw[45] ;
 wire \top_I.branch[13].l_um_iw[46] ;
 wire \top_I.branch[13].l_um_iw[47] ;
 wire \top_I.branch[13].l_um_iw[48] ;
 wire \top_I.branch[13].l_um_iw[49] ;
 wire \top_I.branch[13].l_um_iw[4] ;
 wire \top_I.branch[13].l_um_iw[50] ;
 wire \top_I.branch[13].l_um_iw[51] ;
 wire \top_I.branch[13].l_um_iw[52] ;
 wire \top_I.branch[13].l_um_iw[53] ;
 wire \top_I.branch[13].l_um_iw[54] ;
 wire \top_I.branch[13].l_um_iw[55] ;
 wire \top_I.branch[13].l_um_iw[56] ;
 wire \top_I.branch[13].l_um_iw[57] ;
 wire \top_I.branch[13].l_um_iw[58] ;
 wire \top_I.branch[13].l_um_iw[59] ;
 wire \top_I.branch[13].l_um_iw[5] ;
 wire \top_I.branch[13].l_um_iw[60] ;
 wire \top_I.branch[13].l_um_iw[61] ;
 wire \top_I.branch[13].l_um_iw[62] ;
 wire \top_I.branch[13].l_um_iw[63] ;
 wire \top_I.branch[13].l_um_iw[64] ;
 wire \top_I.branch[13].l_um_iw[65] ;
 wire \top_I.branch[13].l_um_iw[66] ;
 wire \top_I.branch[13].l_um_iw[67] ;
 wire \top_I.branch[13].l_um_iw[68] ;
 wire \top_I.branch[13].l_um_iw[69] ;
 wire \top_I.branch[13].l_um_iw[6] ;
 wire \top_I.branch[13].l_um_iw[70] ;
 wire \top_I.branch[13].l_um_iw[71] ;
 wire \top_I.branch[13].l_um_iw[72] ;
 wire \top_I.branch[13].l_um_iw[73] ;
 wire \top_I.branch[13].l_um_iw[74] ;
 wire \top_I.branch[13].l_um_iw[75] ;
 wire \top_I.branch[13].l_um_iw[76] ;
 wire \top_I.branch[13].l_um_iw[77] ;
 wire \top_I.branch[13].l_um_iw[78] ;
 wire \top_I.branch[13].l_um_iw[79] ;
 wire \top_I.branch[13].l_um_iw[7] ;
 wire \top_I.branch[13].l_um_iw[80] ;
 wire \top_I.branch[13].l_um_iw[81] ;
 wire \top_I.branch[13].l_um_iw[82] ;
 wire \top_I.branch[13].l_um_iw[83] ;
 wire \top_I.branch[13].l_um_iw[84] ;
 wire \top_I.branch[13].l_um_iw[85] ;
 wire \top_I.branch[13].l_um_iw[86] ;
 wire \top_I.branch[13].l_um_iw[87] ;
 wire \top_I.branch[13].l_um_iw[88] ;
 wire \top_I.branch[13].l_um_iw[89] ;
 wire \top_I.branch[13].l_um_iw[8] ;
 wire \top_I.branch[13].l_um_iw[90] ;
 wire \top_I.branch[13].l_um_iw[91] ;
 wire \top_I.branch[13].l_um_iw[92] ;
 wire \top_I.branch[13].l_um_iw[93] ;
 wire \top_I.branch[13].l_um_iw[94] ;
 wire \top_I.branch[13].l_um_iw[95] ;
 wire \top_I.branch[13].l_um_iw[96] ;
 wire \top_I.branch[13].l_um_iw[97] ;
 wire \top_I.branch[13].l_um_iw[98] ;
 wire \top_I.branch[13].l_um_iw[99] ;
 wire \top_I.branch[13].l_um_iw[9] ;
 wire \top_I.branch[13].l_um_k_zero[0] ;
 wire \top_I.branch[13].l_um_k_zero[10] ;
 wire \top_I.branch[13].l_um_k_zero[11] ;
 wire \top_I.branch[13].l_um_k_zero[12] ;
 wire \top_I.branch[13].l_um_k_zero[13] ;
 wire \top_I.branch[13].l_um_k_zero[14] ;
 wire \top_I.branch[13].l_um_k_zero[15] ;
 wire \top_I.branch[13].l_um_k_zero[1] ;
 wire \top_I.branch[13].l_um_k_zero[2] ;
 wire \top_I.branch[13].l_um_k_zero[3] ;
 wire \top_I.branch[13].l_um_k_zero[4] ;
 wire \top_I.branch[13].l_um_k_zero[5] ;
 wire \top_I.branch[13].l_um_k_zero[6] ;
 wire \top_I.branch[13].l_um_k_zero[7] ;
 wire \top_I.branch[13].l_um_k_zero[8] ;
 wire \top_I.branch[13].l_um_k_zero[9] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[14].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[14].l_k_one ;
 wire \top_I.branch[14].l_k_zero ;
 wire \top_I.branch[14].l_um_ena[0] ;
 wire \top_I.branch[14].l_um_ena[10] ;
 wire \top_I.branch[14].l_um_ena[11] ;
 wire \top_I.branch[14].l_um_ena[12] ;
 wire \top_I.branch[14].l_um_ena[13] ;
 wire \top_I.branch[14].l_um_ena[14] ;
 wire \top_I.branch[14].l_um_ena[15] ;
 wire \top_I.branch[14].l_um_ena[1] ;
 wire \top_I.branch[14].l_um_ena[2] ;
 wire \top_I.branch[14].l_um_ena[3] ;
 wire \top_I.branch[14].l_um_ena[4] ;
 wire \top_I.branch[14].l_um_ena[5] ;
 wire \top_I.branch[14].l_um_ena[6] ;
 wire \top_I.branch[14].l_um_ena[7] ;
 wire \top_I.branch[14].l_um_ena[8] ;
 wire \top_I.branch[14].l_um_ena[9] ;
 wire \top_I.branch[14].l_um_iw[0] ;
 wire \top_I.branch[14].l_um_iw[100] ;
 wire \top_I.branch[14].l_um_iw[101] ;
 wire \top_I.branch[14].l_um_iw[102] ;
 wire \top_I.branch[14].l_um_iw[103] ;
 wire \top_I.branch[14].l_um_iw[104] ;
 wire \top_I.branch[14].l_um_iw[105] ;
 wire \top_I.branch[14].l_um_iw[106] ;
 wire \top_I.branch[14].l_um_iw[107] ;
 wire \top_I.branch[14].l_um_iw[108] ;
 wire \top_I.branch[14].l_um_iw[109] ;
 wire \top_I.branch[14].l_um_iw[10] ;
 wire \top_I.branch[14].l_um_iw[110] ;
 wire \top_I.branch[14].l_um_iw[111] ;
 wire \top_I.branch[14].l_um_iw[112] ;
 wire \top_I.branch[14].l_um_iw[113] ;
 wire \top_I.branch[14].l_um_iw[114] ;
 wire \top_I.branch[14].l_um_iw[115] ;
 wire \top_I.branch[14].l_um_iw[116] ;
 wire \top_I.branch[14].l_um_iw[117] ;
 wire \top_I.branch[14].l_um_iw[118] ;
 wire \top_I.branch[14].l_um_iw[119] ;
 wire \top_I.branch[14].l_um_iw[11] ;
 wire \top_I.branch[14].l_um_iw[120] ;
 wire \top_I.branch[14].l_um_iw[121] ;
 wire \top_I.branch[14].l_um_iw[122] ;
 wire \top_I.branch[14].l_um_iw[123] ;
 wire \top_I.branch[14].l_um_iw[124] ;
 wire \top_I.branch[14].l_um_iw[125] ;
 wire \top_I.branch[14].l_um_iw[126] ;
 wire \top_I.branch[14].l_um_iw[127] ;
 wire \top_I.branch[14].l_um_iw[128] ;
 wire \top_I.branch[14].l_um_iw[129] ;
 wire \top_I.branch[14].l_um_iw[12] ;
 wire \top_I.branch[14].l_um_iw[130] ;
 wire \top_I.branch[14].l_um_iw[131] ;
 wire \top_I.branch[14].l_um_iw[132] ;
 wire \top_I.branch[14].l_um_iw[133] ;
 wire \top_I.branch[14].l_um_iw[134] ;
 wire \top_I.branch[14].l_um_iw[135] ;
 wire \top_I.branch[14].l_um_iw[136] ;
 wire \top_I.branch[14].l_um_iw[137] ;
 wire \top_I.branch[14].l_um_iw[138] ;
 wire \top_I.branch[14].l_um_iw[139] ;
 wire \top_I.branch[14].l_um_iw[13] ;
 wire \top_I.branch[14].l_um_iw[140] ;
 wire \top_I.branch[14].l_um_iw[141] ;
 wire \top_I.branch[14].l_um_iw[142] ;
 wire \top_I.branch[14].l_um_iw[143] ;
 wire \top_I.branch[14].l_um_iw[144] ;
 wire \top_I.branch[14].l_um_iw[145] ;
 wire \top_I.branch[14].l_um_iw[146] ;
 wire \top_I.branch[14].l_um_iw[147] ;
 wire \top_I.branch[14].l_um_iw[148] ;
 wire \top_I.branch[14].l_um_iw[149] ;
 wire \top_I.branch[14].l_um_iw[14] ;
 wire \top_I.branch[14].l_um_iw[150] ;
 wire \top_I.branch[14].l_um_iw[151] ;
 wire \top_I.branch[14].l_um_iw[152] ;
 wire \top_I.branch[14].l_um_iw[153] ;
 wire \top_I.branch[14].l_um_iw[154] ;
 wire \top_I.branch[14].l_um_iw[155] ;
 wire \top_I.branch[14].l_um_iw[156] ;
 wire \top_I.branch[14].l_um_iw[157] ;
 wire \top_I.branch[14].l_um_iw[158] ;
 wire \top_I.branch[14].l_um_iw[159] ;
 wire \top_I.branch[14].l_um_iw[15] ;
 wire \top_I.branch[14].l_um_iw[160] ;
 wire \top_I.branch[14].l_um_iw[161] ;
 wire \top_I.branch[14].l_um_iw[162] ;
 wire \top_I.branch[14].l_um_iw[163] ;
 wire \top_I.branch[14].l_um_iw[164] ;
 wire \top_I.branch[14].l_um_iw[165] ;
 wire \top_I.branch[14].l_um_iw[166] ;
 wire \top_I.branch[14].l_um_iw[167] ;
 wire \top_I.branch[14].l_um_iw[168] ;
 wire \top_I.branch[14].l_um_iw[169] ;
 wire \top_I.branch[14].l_um_iw[16] ;
 wire \top_I.branch[14].l_um_iw[170] ;
 wire \top_I.branch[14].l_um_iw[171] ;
 wire \top_I.branch[14].l_um_iw[172] ;
 wire \top_I.branch[14].l_um_iw[173] ;
 wire \top_I.branch[14].l_um_iw[174] ;
 wire \top_I.branch[14].l_um_iw[175] ;
 wire \top_I.branch[14].l_um_iw[176] ;
 wire \top_I.branch[14].l_um_iw[177] ;
 wire \top_I.branch[14].l_um_iw[178] ;
 wire \top_I.branch[14].l_um_iw[179] ;
 wire \top_I.branch[14].l_um_iw[17] ;
 wire \top_I.branch[14].l_um_iw[180] ;
 wire \top_I.branch[14].l_um_iw[181] ;
 wire \top_I.branch[14].l_um_iw[182] ;
 wire \top_I.branch[14].l_um_iw[183] ;
 wire \top_I.branch[14].l_um_iw[184] ;
 wire \top_I.branch[14].l_um_iw[185] ;
 wire \top_I.branch[14].l_um_iw[186] ;
 wire \top_I.branch[14].l_um_iw[187] ;
 wire \top_I.branch[14].l_um_iw[188] ;
 wire \top_I.branch[14].l_um_iw[189] ;
 wire \top_I.branch[14].l_um_iw[18] ;
 wire \top_I.branch[14].l_um_iw[190] ;
 wire \top_I.branch[14].l_um_iw[191] ;
 wire \top_I.branch[14].l_um_iw[192] ;
 wire \top_I.branch[14].l_um_iw[193] ;
 wire \top_I.branch[14].l_um_iw[194] ;
 wire \top_I.branch[14].l_um_iw[195] ;
 wire \top_I.branch[14].l_um_iw[196] ;
 wire \top_I.branch[14].l_um_iw[197] ;
 wire \top_I.branch[14].l_um_iw[198] ;
 wire \top_I.branch[14].l_um_iw[199] ;
 wire \top_I.branch[14].l_um_iw[19] ;
 wire \top_I.branch[14].l_um_iw[1] ;
 wire \top_I.branch[14].l_um_iw[200] ;
 wire \top_I.branch[14].l_um_iw[201] ;
 wire \top_I.branch[14].l_um_iw[202] ;
 wire \top_I.branch[14].l_um_iw[203] ;
 wire \top_I.branch[14].l_um_iw[204] ;
 wire \top_I.branch[14].l_um_iw[205] ;
 wire \top_I.branch[14].l_um_iw[206] ;
 wire \top_I.branch[14].l_um_iw[207] ;
 wire \top_I.branch[14].l_um_iw[208] ;
 wire \top_I.branch[14].l_um_iw[209] ;
 wire \top_I.branch[14].l_um_iw[20] ;
 wire \top_I.branch[14].l_um_iw[210] ;
 wire \top_I.branch[14].l_um_iw[211] ;
 wire \top_I.branch[14].l_um_iw[212] ;
 wire \top_I.branch[14].l_um_iw[213] ;
 wire \top_I.branch[14].l_um_iw[214] ;
 wire \top_I.branch[14].l_um_iw[215] ;
 wire \top_I.branch[14].l_um_iw[216] ;
 wire \top_I.branch[14].l_um_iw[217] ;
 wire \top_I.branch[14].l_um_iw[218] ;
 wire \top_I.branch[14].l_um_iw[219] ;
 wire \top_I.branch[14].l_um_iw[21] ;
 wire \top_I.branch[14].l_um_iw[220] ;
 wire \top_I.branch[14].l_um_iw[221] ;
 wire \top_I.branch[14].l_um_iw[222] ;
 wire \top_I.branch[14].l_um_iw[223] ;
 wire \top_I.branch[14].l_um_iw[224] ;
 wire \top_I.branch[14].l_um_iw[225] ;
 wire \top_I.branch[14].l_um_iw[226] ;
 wire \top_I.branch[14].l_um_iw[227] ;
 wire \top_I.branch[14].l_um_iw[228] ;
 wire \top_I.branch[14].l_um_iw[229] ;
 wire \top_I.branch[14].l_um_iw[22] ;
 wire \top_I.branch[14].l_um_iw[230] ;
 wire \top_I.branch[14].l_um_iw[231] ;
 wire \top_I.branch[14].l_um_iw[232] ;
 wire \top_I.branch[14].l_um_iw[233] ;
 wire \top_I.branch[14].l_um_iw[234] ;
 wire \top_I.branch[14].l_um_iw[235] ;
 wire \top_I.branch[14].l_um_iw[236] ;
 wire \top_I.branch[14].l_um_iw[237] ;
 wire \top_I.branch[14].l_um_iw[238] ;
 wire \top_I.branch[14].l_um_iw[239] ;
 wire \top_I.branch[14].l_um_iw[23] ;
 wire \top_I.branch[14].l_um_iw[240] ;
 wire \top_I.branch[14].l_um_iw[241] ;
 wire \top_I.branch[14].l_um_iw[242] ;
 wire \top_I.branch[14].l_um_iw[243] ;
 wire \top_I.branch[14].l_um_iw[244] ;
 wire \top_I.branch[14].l_um_iw[245] ;
 wire \top_I.branch[14].l_um_iw[246] ;
 wire \top_I.branch[14].l_um_iw[247] ;
 wire \top_I.branch[14].l_um_iw[248] ;
 wire \top_I.branch[14].l_um_iw[249] ;
 wire \top_I.branch[14].l_um_iw[24] ;
 wire \top_I.branch[14].l_um_iw[250] ;
 wire \top_I.branch[14].l_um_iw[251] ;
 wire \top_I.branch[14].l_um_iw[252] ;
 wire \top_I.branch[14].l_um_iw[253] ;
 wire \top_I.branch[14].l_um_iw[254] ;
 wire \top_I.branch[14].l_um_iw[255] ;
 wire \top_I.branch[14].l_um_iw[256] ;
 wire \top_I.branch[14].l_um_iw[257] ;
 wire \top_I.branch[14].l_um_iw[258] ;
 wire \top_I.branch[14].l_um_iw[259] ;
 wire \top_I.branch[14].l_um_iw[25] ;
 wire \top_I.branch[14].l_um_iw[260] ;
 wire \top_I.branch[14].l_um_iw[261] ;
 wire \top_I.branch[14].l_um_iw[262] ;
 wire \top_I.branch[14].l_um_iw[263] ;
 wire \top_I.branch[14].l_um_iw[264] ;
 wire \top_I.branch[14].l_um_iw[265] ;
 wire \top_I.branch[14].l_um_iw[266] ;
 wire \top_I.branch[14].l_um_iw[267] ;
 wire \top_I.branch[14].l_um_iw[268] ;
 wire \top_I.branch[14].l_um_iw[269] ;
 wire \top_I.branch[14].l_um_iw[26] ;
 wire \top_I.branch[14].l_um_iw[270] ;
 wire \top_I.branch[14].l_um_iw[271] ;
 wire \top_I.branch[14].l_um_iw[272] ;
 wire \top_I.branch[14].l_um_iw[273] ;
 wire \top_I.branch[14].l_um_iw[274] ;
 wire \top_I.branch[14].l_um_iw[275] ;
 wire \top_I.branch[14].l_um_iw[276] ;
 wire \top_I.branch[14].l_um_iw[277] ;
 wire \top_I.branch[14].l_um_iw[278] ;
 wire \top_I.branch[14].l_um_iw[279] ;
 wire \top_I.branch[14].l_um_iw[27] ;
 wire \top_I.branch[14].l_um_iw[280] ;
 wire \top_I.branch[14].l_um_iw[281] ;
 wire \top_I.branch[14].l_um_iw[282] ;
 wire \top_I.branch[14].l_um_iw[283] ;
 wire \top_I.branch[14].l_um_iw[284] ;
 wire \top_I.branch[14].l_um_iw[285] ;
 wire \top_I.branch[14].l_um_iw[286] ;
 wire \top_I.branch[14].l_um_iw[287] ;
 wire \top_I.branch[14].l_um_iw[28] ;
 wire \top_I.branch[14].l_um_iw[29] ;
 wire \top_I.branch[14].l_um_iw[2] ;
 wire \top_I.branch[14].l_um_iw[30] ;
 wire \top_I.branch[14].l_um_iw[31] ;
 wire \top_I.branch[14].l_um_iw[32] ;
 wire \top_I.branch[14].l_um_iw[33] ;
 wire \top_I.branch[14].l_um_iw[34] ;
 wire \top_I.branch[14].l_um_iw[35] ;
 wire \top_I.branch[14].l_um_iw[36] ;
 wire \top_I.branch[14].l_um_iw[37] ;
 wire \top_I.branch[14].l_um_iw[38] ;
 wire \top_I.branch[14].l_um_iw[39] ;
 wire \top_I.branch[14].l_um_iw[3] ;
 wire \top_I.branch[14].l_um_iw[40] ;
 wire \top_I.branch[14].l_um_iw[41] ;
 wire \top_I.branch[14].l_um_iw[42] ;
 wire \top_I.branch[14].l_um_iw[43] ;
 wire \top_I.branch[14].l_um_iw[44] ;
 wire \top_I.branch[14].l_um_iw[45] ;
 wire \top_I.branch[14].l_um_iw[46] ;
 wire \top_I.branch[14].l_um_iw[47] ;
 wire \top_I.branch[14].l_um_iw[48] ;
 wire \top_I.branch[14].l_um_iw[49] ;
 wire \top_I.branch[14].l_um_iw[4] ;
 wire \top_I.branch[14].l_um_iw[50] ;
 wire \top_I.branch[14].l_um_iw[51] ;
 wire \top_I.branch[14].l_um_iw[52] ;
 wire \top_I.branch[14].l_um_iw[53] ;
 wire \top_I.branch[14].l_um_iw[54] ;
 wire \top_I.branch[14].l_um_iw[55] ;
 wire \top_I.branch[14].l_um_iw[56] ;
 wire \top_I.branch[14].l_um_iw[57] ;
 wire \top_I.branch[14].l_um_iw[58] ;
 wire \top_I.branch[14].l_um_iw[59] ;
 wire \top_I.branch[14].l_um_iw[5] ;
 wire \top_I.branch[14].l_um_iw[60] ;
 wire \top_I.branch[14].l_um_iw[61] ;
 wire \top_I.branch[14].l_um_iw[62] ;
 wire \top_I.branch[14].l_um_iw[63] ;
 wire \top_I.branch[14].l_um_iw[64] ;
 wire \top_I.branch[14].l_um_iw[65] ;
 wire \top_I.branch[14].l_um_iw[66] ;
 wire \top_I.branch[14].l_um_iw[67] ;
 wire \top_I.branch[14].l_um_iw[68] ;
 wire \top_I.branch[14].l_um_iw[69] ;
 wire \top_I.branch[14].l_um_iw[6] ;
 wire \top_I.branch[14].l_um_iw[70] ;
 wire \top_I.branch[14].l_um_iw[71] ;
 wire \top_I.branch[14].l_um_iw[72] ;
 wire \top_I.branch[14].l_um_iw[73] ;
 wire \top_I.branch[14].l_um_iw[74] ;
 wire \top_I.branch[14].l_um_iw[75] ;
 wire \top_I.branch[14].l_um_iw[76] ;
 wire \top_I.branch[14].l_um_iw[77] ;
 wire \top_I.branch[14].l_um_iw[78] ;
 wire \top_I.branch[14].l_um_iw[79] ;
 wire \top_I.branch[14].l_um_iw[7] ;
 wire \top_I.branch[14].l_um_iw[80] ;
 wire \top_I.branch[14].l_um_iw[81] ;
 wire \top_I.branch[14].l_um_iw[82] ;
 wire \top_I.branch[14].l_um_iw[83] ;
 wire \top_I.branch[14].l_um_iw[84] ;
 wire \top_I.branch[14].l_um_iw[85] ;
 wire \top_I.branch[14].l_um_iw[86] ;
 wire \top_I.branch[14].l_um_iw[87] ;
 wire \top_I.branch[14].l_um_iw[88] ;
 wire \top_I.branch[14].l_um_iw[89] ;
 wire \top_I.branch[14].l_um_iw[8] ;
 wire \top_I.branch[14].l_um_iw[90] ;
 wire \top_I.branch[14].l_um_iw[91] ;
 wire \top_I.branch[14].l_um_iw[92] ;
 wire \top_I.branch[14].l_um_iw[93] ;
 wire \top_I.branch[14].l_um_iw[94] ;
 wire \top_I.branch[14].l_um_iw[95] ;
 wire \top_I.branch[14].l_um_iw[96] ;
 wire \top_I.branch[14].l_um_iw[97] ;
 wire \top_I.branch[14].l_um_iw[98] ;
 wire \top_I.branch[14].l_um_iw[99] ;
 wire \top_I.branch[14].l_um_iw[9] ;
 wire \top_I.branch[14].l_um_k_zero[0] ;
 wire \top_I.branch[14].l_um_k_zero[10] ;
 wire \top_I.branch[14].l_um_k_zero[11] ;
 wire \top_I.branch[14].l_um_k_zero[12] ;
 wire \top_I.branch[14].l_um_k_zero[13] ;
 wire \top_I.branch[14].l_um_k_zero[14] ;
 wire \top_I.branch[14].l_um_k_zero[15] ;
 wire \top_I.branch[14].l_um_k_zero[1] ;
 wire \top_I.branch[14].l_um_k_zero[2] ;
 wire \top_I.branch[14].l_um_k_zero[3] ;
 wire \top_I.branch[14].l_um_k_zero[4] ;
 wire \top_I.branch[14].l_um_k_zero[5] ;
 wire \top_I.branch[14].l_um_k_zero[6] ;
 wire \top_I.branch[14].l_um_k_zero[7] ;
 wire \top_I.branch[14].l_um_k_zero[8] ;
 wire \top_I.branch[14].l_um_k_zero[9] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[15].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[15].l_k_one ;
 wire \top_I.branch[15].l_k_zero ;
 wire \top_I.branch[15].l_um_ena[0] ;
 wire \top_I.branch[15].l_um_ena[10] ;
 wire \top_I.branch[15].l_um_ena[11] ;
 wire \top_I.branch[15].l_um_ena[12] ;
 wire \top_I.branch[15].l_um_ena[13] ;
 wire \top_I.branch[15].l_um_ena[14] ;
 wire \top_I.branch[15].l_um_ena[15] ;
 wire \top_I.branch[15].l_um_ena[1] ;
 wire \top_I.branch[15].l_um_ena[2] ;
 wire \top_I.branch[15].l_um_ena[3] ;
 wire \top_I.branch[15].l_um_ena[4] ;
 wire \top_I.branch[15].l_um_ena[5] ;
 wire \top_I.branch[15].l_um_ena[6] ;
 wire \top_I.branch[15].l_um_ena[7] ;
 wire \top_I.branch[15].l_um_ena[8] ;
 wire \top_I.branch[15].l_um_ena[9] ;
 wire \top_I.branch[15].l_um_iw[0] ;
 wire \top_I.branch[15].l_um_iw[100] ;
 wire \top_I.branch[15].l_um_iw[101] ;
 wire \top_I.branch[15].l_um_iw[102] ;
 wire \top_I.branch[15].l_um_iw[103] ;
 wire \top_I.branch[15].l_um_iw[104] ;
 wire \top_I.branch[15].l_um_iw[105] ;
 wire \top_I.branch[15].l_um_iw[106] ;
 wire \top_I.branch[15].l_um_iw[107] ;
 wire \top_I.branch[15].l_um_iw[108] ;
 wire \top_I.branch[15].l_um_iw[109] ;
 wire \top_I.branch[15].l_um_iw[10] ;
 wire \top_I.branch[15].l_um_iw[110] ;
 wire \top_I.branch[15].l_um_iw[111] ;
 wire \top_I.branch[15].l_um_iw[112] ;
 wire \top_I.branch[15].l_um_iw[113] ;
 wire \top_I.branch[15].l_um_iw[114] ;
 wire \top_I.branch[15].l_um_iw[115] ;
 wire \top_I.branch[15].l_um_iw[116] ;
 wire \top_I.branch[15].l_um_iw[117] ;
 wire \top_I.branch[15].l_um_iw[118] ;
 wire \top_I.branch[15].l_um_iw[119] ;
 wire \top_I.branch[15].l_um_iw[11] ;
 wire \top_I.branch[15].l_um_iw[120] ;
 wire \top_I.branch[15].l_um_iw[121] ;
 wire \top_I.branch[15].l_um_iw[122] ;
 wire \top_I.branch[15].l_um_iw[123] ;
 wire \top_I.branch[15].l_um_iw[124] ;
 wire \top_I.branch[15].l_um_iw[125] ;
 wire \top_I.branch[15].l_um_iw[126] ;
 wire \top_I.branch[15].l_um_iw[127] ;
 wire \top_I.branch[15].l_um_iw[128] ;
 wire \top_I.branch[15].l_um_iw[129] ;
 wire \top_I.branch[15].l_um_iw[12] ;
 wire \top_I.branch[15].l_um_iw[130] ;
 wire \top_I.branch[15].l_um_iw[131] ;
 wire \top_I.branch[15].l_um_iw[132] ;
 wire \top_I.branch[15].l_um_iw[133] ;
 wire \top_I.branch[15].l_um_iw[134] ;
 wire \top_I.branch[15].l_um_iw[135] ;
 wire \top_I.branch[15].l_um_iw[136] ;
 wire \top_I.branch[15].l_um_iw[137] ;
 wire \top_I.branch[15].l_um_iw[138] ;
 wire \top_I.branch[15].l_um_iw[139] ;
 wire \top_I.branch[15].l_um_iw[13] ;
 wire \top_I.branch[15].l_um_iw[140] ;
 wire \top_I.branch[15].l_um_iw[141] ;
 wire \top_I.branch[15].l_um_iw[142] ;
 wire \top_I.branch[15].l_um_iw[143] ;
 wire \top_I.branch[15].l_um_iw[144] ;
 wire \top_I.branch[15].l_um_iw[145] ;
 wire \top_I.branch[15].l_um_iw[146] ;
 wire \top_I.branch[15].l_um_iw[147] ;
 wire \top_I.branch[15].l_um_iw[148] ;
 wire \top_I.branch[15].l_um_iw[149] ;
 wire \top_I.branch[15].l_um_iw[14] ;
 wire \top_I.branch[15].l_um_iw[150] ;
 wire \top_I.branch[15].l_um_iw[151] ;
 wire \top_I.branch[15].l_um_iw[152] ;
 wire \top_I.branch[15].l_um_iw[153] ;
 wire \top_I.branch[15].l_um_iw[154] ;
 wire \top_I.branch[15].l_um_iw[155] ;
 wire \top_I.branch[15].l_um_iw[156] ;
 wire \top_I.branch[15].l_um_iw[157] ;
 wire \top_I.branch[15].l_um_iw[158] ;
 wire \top_I.branch[15].l_um_iw[159] ;
 wire \top_I.branch[15].l_um_iw[15] ;
 wire \top_I.branch[15].l_um_iw[160] ;
 wire \top_I.branch[15].l_um_iw[161] ;
 wire \top_I.branch[15].l_um_iw[162] ;
 wire \top_I.branch[15].l_um_iw[163] ;
 wire \top_I.branch[15].l_um_iw[164] ;
 wire \top_I.branch[15].l_um_iw[165] ;
 wire \top_I.branch[15].l_um_iw[166] ;
 wire \top_I.branch[15].l_um_iw[167] ;
 wire \top_I.branch[15].l_um_iw[168] ;
 wire \top_I.branch[15].l_um_iw[169] ;
 wire \top_I.branch[15].l_um_iw[16] ;
 wire \top_I.branch[15].l_um_iw[170] ;
 wire \top_I.branch[15].l_um_iw[171] ;
 wire \top_I.branch[15].l_um_iw[172] ;
 wire \top_I.branch[15].l_um_iw[173] ;
 wire \top_I.branch[15].l_um_iw[174] ;
 wire \top_I.branch[15].l_um_iw[175] ;
 wire \top_I.branch[15].l_um_iw[176] ;
 wire \top_I.branch[15].l_um_iw[177] ;
 wire \top_I.branch[15].l_um_iw[178] ;
 wire \top_I.branch[15].l_um_iw[179] ;
 wire \top_I.branch[15].l_um_iw[17] ;
 wire \top_I.branch[15].l_um_iw[180] ;
 wire \top_I.branch[15].l_um_iw[181] ;
 wire \top_I.branch[15].l_um_iw[182] ;
 wire \top_I.branch[15].l_um_iw[183] ;
 wire \top_I.branch[15].l_um_iw[184] ;
 wire \top_I.branch[15].l_um_iw[185] ;
 wire \top_I.branch[15].l_um_iw[186] ;
 wire \top_I.branch[15].l_um_iw[187] ;
 wire \top_I.branch[15].l_um_iw[188] ;
 wire \top_I.branch[15].l_um_iw[189] ;
 wire \top_I.branch[15].l_um_iw[18] ;
 wire \top_I.branch[15].l_um_iw[190] ;
 wire \top_I.branch[15].l_um_iw[191] ;
 wire \top_I.branch[15].l_um_iw[192] ;
 wire \top_I.branch[15].l_um_iw[193] ;
 wire \top_I.branch[15].l_um_iw[194] ;
 wire \top_I.branch[15].l_um_iw[195] ;
 wire \top_I.branch[15].l_um_iw[196] ;
 wire \top_I.branch[15].l_um_iw[197] ;
 wire \top_I.branch[15].l_um_iw[198] ;
 wire \top_I.branch[15].l_um_iw[199] ;
 wire \top_I.branch[15].l_um_iw[19] ;
 wire \top_I.branch[15].l_um_iw[1] ;
 wire \top_I.branch[15].l_um_iw[200] ;
 wire \top_I.branch[15].l_um_iw[201] ;
 wire \top_I.branch[15].l_um_iw[202] ;
 wire \top_I.branch[15].l_um_iw[203] ;
 wire \top_I.branch[15].l_um_iw[204] ;
 wire \top_I.branch[15].l_um_iw[205] ;
 wire \top_I.branch[15].l_um_iw[206] ;
 wire \top_I.branch[15].l_um_iw[207] ;
 wire \top_I.branch[15].l_um_iw[208] ;
 wire \top_I.branch[15].l_um_iw[209] ;
 wire \top_I.branch[15].l_um_iw[20] ;
 wire \top_I.branch[15].l_um_iw[210] ;
 wire \top_I.branch[15].l_um_iw[211] ;
 wire \top_I.branch[15].l_um_iw[212] ;
 wire \top_I.branch[15].l_um_iw[213] ;
 wire \top_I.branch[15].l_um_iw[214] ;
 wire \top_I.branch[15].l_um_iw[215] ;
 wire \top_I.branch[15].l_um_iw[216] ;
 wire \top_I.branch[15].l_um_iw[217] ;
 wire \top_I.branch[15].l_um_iw[218] ;
 wire \top_I.branch[15].l_um_iw[219] ;
 wire \top_I.branch[15].l_um_iw[21] ;
 wire \top_I.branch[15].l_um_iw[220] ;
 wire \top_I.branch[15].l_um_iw[221] ;
 wire \top_I.branch[15].l_um_iw[222] ;
 wire \top_I.branch[15].l_um_iw[223] ;
 wire \top_I.branch[15].l_um_iw[224] ;
 wire \top_I.branch[15].l_um_iw[225] ;
 wire \top_I.branch[15].l_um_iw[226] ;
 wire \top_I.branch[15].l_um_iw[227] ;
 wire \top_I.branch[15].l_um_iw[228] ;
 wire \top_I.branch[15].l_um_iw[229] ;
 wire \top_I.branch[15].l_um_iw[22] ;
 wire \top_I.branch[15].l_um_iw[230] ;
 wire \top_I.branch[15].l_um_iw[231] ;
 wire \top_I.branch[15].l_um_iw[232] ;
 wire \top_I.branch[15].l_um_iw[233] ;
 wire \top_I.branch[15].l_um_iw[234] ;
 wire \top_I.branch[15].l_um_iw[235] ;
 wire \top_I.branch[15].l_um_iw[236] ;
 wire \top_I.branch[15].l_um_iw[237] ;
 wire \top_I.branch[15].l_um_iw[238] ;
 wire \top_I.branch[15].l_um_iw[239] ;
 wire \top_I.branch[15].l_um_iw[23] ;
 wire \top_I.branch[15].l_um_iw[240] ;
 wire \top_I.branch[15].l_um_iw[241] ;
 wire \top_I.branch[15].l_um_iw[242] ;
 wire \top_I.branch[15].l_um_iw[243] ;
 wire \top_I.branch[15].l_um_iw[244] ;
 wire \top_I.branch[15].l_um_iw[245] ;
 wire \top_I.branch[15].l_um_iw[246] ;
 wire \top_I.branch[15].l_um_iw[247] ;
 wire \top_I.branch[15].l_um_iw[248] ;
 wire \top_I.branch[15].l_um_iw[249] ;
 wire \top_I.branch[15].l_um_iw[24] ;
 wire \top_I.branch[15].l_um_iw[250] ;
 wire \top_I.branch[15].l_um_iw[251] ;
 wire \top_I.branch[15].l_um_iw[252] ;
 wire \top_I.branch[15].l_um_iw[253] ;
 wire \top_I.branch[15].l_um_iw[254] ;
 wire \top_I.branch[15].l_um_iw[255] ;
 wire \top_I.branch[15].l_um_iw[256] ;
 wire \top_I.branch[15].l_um_iw[257] ;
 wire \top_I.branch[15].l_um_iw[258] ;
 wire \top_I.branch[15].l_um_iw[259] ;
 wire \top_I.branch[15].l_um_iw[25] ;
 wire \top_I.branch[15].l_um_iw[260] ;
 wire \top_I.branch[15].l_um_iw[261] ;
 wire \top_I.branch[15].l_um_iw[262] ;
 wire \top_I.branch[15].l_um_iw[263] ;
 wire \top_I.branch[15].l_um_iw[264] ;
 wire \top_I.branch[15].l_um_iw[265] ;
 wire \top_I.branch[15].l_um_iw[266] ;
 wire \top_I.branch[15].l_um_iw[267] ;
 wire \top_I.branch[15].l_um_iw[268] ;
 wire \top_I.branch[15].l_um_iw[269] ;
 wire \top_I.branch[15].l_um_iw[26] ;
 wire \top_I.branch[15].l_um_iw[270] ;
 wire \top_I.branch[15].l_um_iw[271] ;
 wire \top_I.branch[15].l_um_iw[272] ;
 wire \top_I.branch[15].l_um_iw[273] ;
 wire \top_I.branch[15].l_um_iw[274] ;
 wire \top_I.branch[15].l_um_iw[275] ;
 wire \top_I.branch[15].l_um_iw[276] ;
 wire \top_I.branch[15].l_um_iw[277] ;
 wire \top_I.branch[15].l_um_iw[278] ;
 wire \top_I.branch[15].l_um_iw[279] ;
 wire \top_I.branch[15].l_um_iw[27] ;
 wire \top_I.branch[15].l_um_iw[280] ;
 wire \top_I.branch[15].l_um_iw[281] ;
 wire \top_I.branch[15].l_um_iw[282] ;
 wire \top_I.branch[15].l_um_iw[283] ;
 wire \top_I.branch[15].l_um_iw[284] ;
 wire \top_I.branch[15].l_um_iw[285] ;
 wire \top_I.branch[15].l_um_iw[286] ;
 wire \top_I.branch[15].l_um_iw[287] ;
 wire \top_I.branch[15].l_um_iw[28] ;
 wire \top_I.branch[15].l_um_iw[29] ;
 wire \top_I.branch[15].l_um_iw[2] ;
 wire \top_I.branch[15].l_um_iw[30] ;
 wire \top_I.branch[15].l_um_iw[31] ;
 wire \top_I.branch[15].l_um_iw[32] ;
 wire \top_I.branch[15].l_um_iw[33] ;
 wire \top_I.branch[15].l_um_iw[34] ;
 wire \top_I.branch[15].l_um_iw[35] ;
 wire \top_I.branch[15].l_um_iw[36] ;
 wire \top_I.branch[15].l_um_iw[37] ;
 wire \top_I.branch[15].l_um_iw[38] ;
 wire \top_I.branch[15].l_um_iw[39] ;
 wire \top_I.branch[15].l_um_iw[3] ;
 wire \top_I.branch[15].l_um_iw[40] ;
 wire \top_I.branch[15].l_um_iw[41] ;
 wire \top_I.branch[15].l_um_iw[42] ;
 wire \top_I.branch[15].l_um_iw[43] ;
 wire \top_I.branch[15].l_um_iw[44] ;
 wire \top_I.branch[15].l_um_iw[45] ;
 wire \top_I.branch[15].l_um_iw[46] ;
 wire \top_I.branch[15].l_um_iw[47] ;
 wire \top_I.branch[15].l_um_iw[48] ;
 wire \top_I.branch[15].l_um_iw[49] ;
 wire \top_I.branch[15].l_um_iw[4] ;
 wire \top_I.branch[15].l_um_iw[50] ;
 wire \top_I.branch[15].l_um_iw[51] ;
 wire \top_I.branch[15].l_um_iw[52] ;
 wire \top_I.branch[15].l_um_iw[53] ;
 wire \top_I.branch[15].l_um_iw[54] ;
 wire \top_I.branch[15].l_um_iw[55] ;
 wire \top_I.branch[15].l_um_iw[56] ;
 wire \top_I.branch[15].l_um_iw[57] ;
 wire \top_I.branch[15].l_um_iw[58] ;
 wire \top_I.branch[15].l_um_iw[59] ;
 wire \top_I.branch[15].l_um_iw[5] ;
 wire \top_I.branch[15].l_um_iw[60] ;
 wire \top_I.branch[15].l_um_iw[61] ;
 wire \top_I.branch[15].l_um_iw[62] ;
 wire \top_I.branch[15].l_um_iw[63] ;
 wire \top_I.branch[15].l_um_iw[64] ;
 wire \top_I.branch[15].l_um_iw[65] ;
 wire \top_I.branch[15].l_um_iw[66] ;
 wire \top_I.branch[15].l_um_iw[67] ;
 wire \top_I.branch[15].l_um_iw[68] ;
 wire \top_I.branch[15].l_um_iw[69] ;
 wire \top_I.branch[15].l_um_iw[6] ;
 wire \top_I.branch[15].l_um_iw[70] ;
 wire \top_I.branch[15].l_um_iw[71] ;
 wire \top_I.branch[15].l_um_iw[72] ;
 wire \top_I.branch[15].l_um_iw[73] ;
 wire \top_I.branch[15].l_um_iw[74] ;
 wire \top_I.branch[15].l_um_iw[75] ;
 wire \top_I.branch[15].l_um_iw[76] ;
 wire \top_I.branch[15].l_um_iw[77] ;
 wire \top_I.branch[15].l_um_iw[78] ;
 wire \top_I.branch[15].l_um_iw[79] ;
 wire \top_I.branch[15].l_um_iw[7] ;
 wire \top_I.branch[15].l_um_iw[80] ;
 wire \top_I.branch[15].l_um_iw[81] ;
 wire \top_I.branch[15].l_um_iw[82] ;
 wire \top_I.branch[15].l_um_iw[83] ;
 wire \top_I.branch[15].l_um_iw[84] ;
 wire \top_I.branch[15].l_um_iw[85] ;
 wire \top_I.branch[15].l_um_iw[86] ;
 wire \top_I.branch[15].l_um_iw[87] ;
 wire \top_I.branch[15].l_um_iw[88] ;
 wire \top_I.branch[15].l_um_iw[89] ;
 wire \top_I.branch[15].l_um_iw[8] ;
 wire \top_I.branch[15].l_um_iw[90] ;
 wire \top_I.branch[15].l_um_iw[91] ;
 wire \top_I.branch[15].l_um_iw[92] ;
 wire \top_I.branch[15].l_um_iw[93] ;
 wire \top_I.branch[15].l_um_iw[94] ;
 wire \top_I.branch[15].l_um_iw[95] ;
 wire \top_I.branch[15].l_um_iw[96] ;
 wire \top_I.branch[15].l_um_iw[97] ;
 wire \top_I.branch[15].l_um_iw[98] ;
 wire \top_I.branch[15].l_um_iw[99] ;
 wire \top_I.branch[15].l_um_iw[9] ;
 wire \top_I.branch[15].l_um_k_zero[0] ;
 wire \top_I.branch[15].l_um_k_zero[10] ;
 wire \top_I.branch[15].l_um_k_zero[11] ;
 wire \top_I.branch[15].l_um_k_zero[12] ;
 wire \top_I.branch[15].l_um_k_zero[13] ;
 wire \top_I.branch[15].l_um_k_zero[14] ;
 wire \top_I.branch[15].l_um_k_zero[15] ;
 wire \top_I.branch[15].l_um_k_zero[1] ;
 wire \top_I.branch[15].l_um_k_zero[2] ;
 wire \top_I.branch[15].l_um_k_zero[3] ;
 wire \top_I.branch[15].l_um_k_zero[4] ;
 wire \top_I.branch[15].l_um_k_zero[5] ;
 wire \top_I.branch[15].l_um_k_zero[6] ;
 wire \top_I.branch[15].l_um_k_zero[7] ;
 wire \top_I.branch[15].l_um_k_zero[8] ;
 wire \top_I.branch[15].l_um_k_zero[9] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[16].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[16].l_k_one ;
 wire \top_I.branch[16].l_k_zero ;
 wire \top_I.branch[16].l_um_ena[0] ;
 wire \top_I.branch[16].l_um_ena[10] ;
 wire \top_I.branch[16].l_um_ena[11] ;
 wire \top_I.branch[16].l_um_ena[12] ;
 wire \top_I.branch[16].l_um_ena[13] ;
 wire \top_I.branch[16].l_um_ena[14] ;
 wire \top_I.branch[16].l_um_ena[15] ;
 wire \top_I.branch[16].l_um_ena[1] ;
 wire \top_I.branch[16].l_um_ena[2] ;
 wire \top_I.branch[16].l_um_ena[3] ;
 wire \top_I.branch[16].l_um_ena[4] ;
 wire \top_I.branch[16].l_um_ena[5] ;
 wire \top_I.branch[16].l_um_ena[6] ;
 wire \top_I.branch[16].l_um_ena[7] ;
 wire \top_I.branch[16].l_um_ena[8] ;
 wire \top_I.branch[16].l_um_ena[9] ;
 wire \top_I.branch[16].l_um_iw[0] ;
 wire \top_I.branch[16].l_um_iw[100] ;
 wire \top_I.branch[16].l_um_iw[101] ;
 wire \top_I.branch[16].l_um_iw[102] ;
 wire \top_I.branch[16].l_um_iw[103] ;
 wire \top_I.branch[16].l_um_iw[104] ;
 wire \top_I.branch[16].l_um_iw[105] ;
 wire \top_I.branch[16].l_um_iw[106] ;
 wire \top_I.branch[16].l_um_iw[107] ;
 wire \top_I.branch[16].l_um_iw[108] ;
 wire \top_I.branch[16].l_um_iw[109] ;
 wire \top_I.branch[16].l_um_iw[10] ;
 wire \top_I.branch[16].l_um_iw[110] ;
 wire \top_I.branch[16].l_um_iw[111] ;
 wire \top_I.branch[16].l_um_iw[112] ;
 wire \top_I.branch[16].l_um_iw[113] ;
 wire \top_I.branch[16].l_um_iw[114] ;
 wire \top_I.branch[16].l_um_iw[115] ;
 wire \top_I.branch[16].l_um_iw[116] ;
 wire \top_I.branch[16].l_um_iw[117] ;
 wire \top_I.branch[16].l_um_iw[118] ;
 wire \top_I.branch[16].l_um_iw[119] ;
 wire \top_I.branch[16].l_um_iw[11] ;
 wire \top_I.branch[16].l_um_iw[120] ;
 wire \top_I.branch[16].l_um_iw[121] ;
 wire \top_I.branch[16].l_um_iw[122] ;
 wire \top_I.branch[16].l_um_iw[123] ;
 wire \top_I.branch[16].l_um_iw[124] ;
 wire \top_I.branch[16].l_um_iw[125] ;
 wire \top_I.branch[16].l_um_iw[126] ;
 wire \top_I.branch[16].l_um_iw[127] ;
 wire \top_I.branch[16].l_um_iw[128] ;
 wire \top_I.branch[16].l_um_iw[129] ;
 wire \top_I.branch[16].l_um_iw[12] ;
 wire \top_I.branch[16].l_um_iw[130] ;
 wire \top_I.branch[16].l_um_iw[131] ;
 wire \top_I.branch[16].l_um_iw[132] ;
 wire \top_I.branch[16].l_um_iw[133] ;
 wire \top_I.branch[16].l_um_iw[134] ;
 wire \top_I.branch[16].l_um_iw[135] ;
 wire \top_I.branch[16].l_um_iw[136] ;
 wire \top_I.branch[16].l_um_iw[137] ;
 wire \top_I.branch[16].l_um_iw[138] ;
 wire \top_I.branch[16].l_um_iw[139] ;
 wire \top_I.branch[16].l_um_iw[13] ;
 wire \top_I.branch[16].l_um_iw[140] ;
 wire \top_I.branch[16].l_um_iw[141] ;
 wire \top_I.branch[16].l_um_iw[142] ;
 wire \top_I.branch[16].l_um_iw[143] ;
 wire \top_I.branch[16].l_um_iw[144] ;
 wire \top_I.branch[16].l_um_iw[145] ;
 wire \top_I.branch[16].l_um_iw[146] ;
 wire \top_I.branch[16].l_um_iw[147] ;
 wire \top_I.branch[16].l_um_iw[148] ;
 wire \top_I.branch[16].l_um_iw[149] ;
 wire \top_I.branch[16].l_um_iw[14] ;
 wire \top_I.branch[16].l_um_iw[150] ;
 wire \top_I.branch[16].l_um_iw[151] ;
 wire \top_I.branch[16].l_um_iw[152] ;
 wire \top_I.branch[16].l_um_iw[153] ;
 wire \top_I.branch[16].l_um_iw[154] ;
 wire \top_I.branch[16].l_um_iw[155] ;
 wire \top_I.branch[16].l_um_iw[156] ;
 wire \top_I.branch[16].l_um_iw[157] ;
 wire \top_I.branch[16].l_um_iw[158] ;
 wire \top_I.branch[16].l_um_iw[159] ;
 wire \top_I.branch[16].l_um_iw[15] ;
 wire \top_I.branch[16].l_um_iw[160] ;
 wire \top_I.branch[16].l_um_iw[161] ;
 wire \top_I.branch[16].l_um_iw[162] ;
 wire \top_I.branch[16].l_um_iw[163] ;
 wire \top_I.branch[16].l_um_iw[164] ;
 wire \top_I.branch[16].l_um_iw[165] ;
 wire \top_I.branch[16].l_um_iw[166] ;
 wire \top_I.branch[16].l_um_iw[167] ;
 wire \top_I.branch[16].l_um_iw[168] ;
 wire \top_I.branch[16].l_um_iw[169] ;
 wire \top_I.branch[16].l_um_iw[16] ;
 wire \top_I.branch[16].l_um_iw[170] ;
 wire \top_I.branch[16].l_um_iw[171] ;
 wire \top_I.branch[16].l_um_iw[172] ;
 wire \top_I.branch[16].l_um_iw[173] ;
 wire \top_I.branch[16].l_um_iw[174] ;
 wire \top_I.branch[16].l_um_iw[175] ;
 wire \top_I.branch[16].l_um_iw[176] ;
 wire \top_I.branch[16].l_um_iw[177] ;
 wire \top_I.branch[16].l_um_iw[178] ;
 wire \top_I.branch[16].l_um_iw[179] ;
 wire \top_I.branch[16].l_um_iw[17] ;
 wire \top_I.branch[16].l_um_iw[180] ;
 wire \top_I.branch[16].l_um_iw[181] ;
 wire \top_I.branch[16].l_um_iw[182] ;
 wire \top_I.branch[16].l_um_iw[183] ;
 wire \top_I.branch[16].l_um_iw[184] ;
 wire \top_I.branch[16].l_um_iw[185] ;
 wire \top_I.branch[16].l_um_iw[186] ;
 wire \top_I.branch[16].l_um_iw[187] ;
 wire \top_I.branch[16].l_um_iw[188] ;
 wire \top_I.branch[16].l_um_iw[189] ;
 wire \top_I.branch[16].l_um_iw[18] ;
 wire \top_I.branch[16].l_um_iw[190] ;
 wire \top_I.branch[16].l_um_iw[191] ;
 wire \top_I.branch[16].l_um_iw[192] ;
 wire \top_I.branch[16].l_um_iw[193] ;
 wire \top_I.branch[16].l_um_iw[194] ;
 wire \top_I.branch[16].l_um_iw[195] ;
 wire \top_I.branch[16].l_um_iw[196] ;
 wire \top_I.branch[16].l_um_iw[197] ;
 wire \top_I.branch[16].l_um_iw[198] ;
 wire \top_I.branch[16].l_um_iw[199] ;
 wire \top_I.branch[16].l_um_iw[19] ;
 wire \top_I.branch[16].l_um_iw[1] ;
 wire \top_I.branch[16].l_um_iw[200] ;
 wire \top_I.branch[16].l_um_iw[201] ;
 wire \top_I.branch[16].l_um_iw[202] ;
 wire \top_I.branch[16].l_um_iw[203] ;
 wire \top_I.branch[16].l_um_iw[204] ;
 wire \top_I.branch[16].l_um_iw[205] ;
 wire \top_I.branch[16].l_um_iw[206] ;
 wire \top_I.branch[16].l_um_iw[207] ;
 wire \top_I.branch[16].l_um_iw[208] ;
 wire \top_I.branch[16].l_um_iw[209] ;
 wire \top_I.branch[16].l_um_iw[20] ;
 wire \top_I.branch[16].l_um_iw[210] ;
 wire \top_I.branch[16].l_um_iw[211] ;
 wire \top_I.branch[16].l_um_iw[212] ;
 wire \top_I.branch[16].l_um_iw[213] ;
 wire \top_I.branch[16].l_um_iw[214] ;
 wire \top_I.branch[16].l_um_iw[215] ;
 wire \top_I.branch[16].l_um_iw[216] ;
 wire \top_I.branch[16].l_um_iw[217] ;
 wire \top_I.branch[16].l_um_iw[218] ;
 wire \top_I.branch[16].l_um_iw[219] ;
 wire \top_I.branch[16].l_um_iw[21] ;
 wire \top_I.branch[16].l_um_iw[220] ;
 wire \top_I.branch[16].l_um_iw[221] ;
 wire \top_I.branch[16].l_um_iw[222] ;
 wire \top_I.branch[16].l_um_iw[223] ;
 wire \top_I.branch[16].l_um_iw[224] ;
 wire \top_I.branch[16].l_um_iw[225] ;
 wire \top_I.branch[16].l_um_iw[226] ;
 wire \top_I.branch[16].l_um_iw[227] ;
 wire \top_I.branch[16].l_um_iw[228] ;
 wire \top_I.branch[16].l_um_iw[229] ;
 wire \top_I.branch[16].l_um_iw[22] ;
 wire \top_I.branch[16].l_um_iw[230] ;
 wire \top_I.branch[16].l_um_iw[231] ;
 wire \top_I.branch[16].l_um_iw[232] ;
 wire \top_I.branch[16].l_um_iw[233] ;
 wire \top_I.branch[16].l_um_iw[234] ;
 wire \top_I.branch[16].l_um_iw[235] ;
 wire \top_I.branch[16].l_um_iw[236] ;
 wire \top_I.branch[16].l_um_iw[237] ;
 wire \top_I.branch[16].l_um_iw[238] ;
 wire \top_I.branch[16].l_um_iw[239] ;
 wire \top_I.branch[16].l_um_iw[23] ;
 wire \top_I.branch[16].l_um_iw[240] ;
 wire \top_I.branch[16].l_um_iw[241] ;
 wire \top_I.branch[16].l_um_iw[242] ;
 wire \top_I.branch[16].l_um_iw[243] ;
 wire \top_I.branch[16].l_um_iw[244] ;
 wire \top_I.branch[16].l_um_iw[245] ;
 wire \top_I.branch[16].l_um_iw[246] ;
 wire \top_I.branch[16].l_um_iw[247] ;
 wire \top_I.branch[16].l_um_iw[248] ;
 wire \top_I.branch[16].l_um_iw[249] ;
 wire \top_I.branch[16].l_um_iw[24] ;
 wire \top_I.branch[16].l_um_iw[250] ;
 wire \top_I.branch[16].l_um_iw[251] ;
 wire \top_I.branch[16].l_um_iw[252] ;
 wire \top_I.branch[16].l_um_iw[253] ;
 wire \top_I.branch[16].l_um_iw[254] ;
 wire \top_I.branch[16].l_um_iw[255] ;
 wire \top_I.branch[16].l_um_iw[256] ;
 wire \top_I.branch[16].l_um_iw[257] ;
 wire \top_I.branch[16].l_um_iw[258] ;
 wire \top_I.branch[16].l_um_iw[259] ;
 wire \top_I.branch[16].l_um_iw[25] ;
 wire \top_I.branch[16].l_um_iw[260] ;
 wire \top_I.branch[16].l_um_iw[261] ;
 wire \top_I.branch[16].l_um_iw[262] ;
 wire \top_I.branch[16].l_um_iw[263] ;
 wire \top_I.branch[16].l_um_iw[264] ;
 wire \top_I.branch[16].l_um_iw[265] ;
 wire \top_I.branch[16].l_um_iw[266] ;
 wire \top_I.branch[16].l_um_iw[267] ;
 wire \top_I.branch[16].l_um_iw[268] ;
 wire \top_I.branch[16].l_um_iw[269] ;
 wire \top_I.branch[16].l_um_iw[26] ;
 wire \top_I.branch[16].l_um_iw[270] ;
 wire \top_I.branch[16].l_um_iw[271] ;
 wire \top_I.branch[16].l_um_iw[272] ;
 wire \top_I.branch[16].l_um_iw[273] ;
 wire \top_I.branch[16].l_um_iw[274] ;
 wire \top_I.branch[16].l_um_iw[275] ;
 wire \top_I.branch[16].l_um_iw[276] ;
 wire \top_I.branch[16].l_um_iw[277] ;
 wire \top_I.branch[16].l_um_iw[278] ;
 wire \top_I.branch[16].l_um_iw[279] ;
 wire \top_I.branch[16].l_um_iw[27] ;
 wire \top_I.branch[16].l_um_iw[280] ;
 wire \top_I.branch[16].l_um_iw[281] ;
 wire \top_I.branch[16].l_um_iw[282] ;
 wire \top_I.branch[16].l_um_iw[283] ;
 wire \top_I.branch[16].l_um_iw[284] ;
 wire \top_I.branch[16].l_um_iw[285] ;
 wire \top_I.branch[16].l_um_iw[286] ;
 wire \top_I.branch[16].l_um_iw[287] ;
 wire \top_I.branch[16].l_um_iw[28] ;
 wire \top_I.branch[16].l_um_iw[29] ;
 wire \top_I.branch[16].l_um_iw[2] ;
 wire \top_I.branch[16].l_um_iw[30] ;
 wire \top_I.branch[16].l_um_iw[31] ;
 wire \top_I.branch[16].l_um_iw[32] ;
 wire \top_I.branch[16].l_um_iw[33] ;
 wire \top_I.branch[16].l_um_iw[34] ;
 wire \top_I.branch[16].l_um_iw[35] ;
 wire \top_I.branch[16].l_um_iw[36] ;
 wire \top_I.branch[16].l_um_iw[37] ;
 wire \top_I.branch[16].l_um_iw[38] ;
 wire \top_I.branch[16].l_um_iw[39] ;
 wire \top_I.branch[16].l_um_iw[3] ;
 wire \top_I.branch[16].l_um_iw[40] ;
 wire \top_I.branch[16].l_um_iw[41] ;
 wire \top_I.branch[16].l_um_iw[42] ;
 wire \top_I.branch[16].l_um_iw[43] ;
 wire \top_I.branch[16].l_um_iw[44] ;
 wire \top_I.branch[16].l_um_iw[45] ;
 wire \top_I.branch[16].l_um_iw[46] ;
 wire \top_I.branch[16].l_um_iw[47] ;
 wire \top_I.branch[16].l_um_iw[48] ;
 wire \top_I.branch[16].l_um_iw[49] ;
 wire \top_I.branch[16].l_um_iw[4] ;
 wire \top_I.branch[16].l_um_iw[50] ;
 wire \top_I.branch[16].l_um_iw[51] ;
 wire \top_I.branch[16].l_um_iw[52] ;
 wire \top_I.branch[16].l_um_iw[53] ;
 wire \top_I.branch[16].l_um_iw[54] ;
 wire \top_I.branch[16].l_um_iw[55] ;
 wire \top_I.branch[16].l_um_iw[56] ;
 wire \top_I.branch[16].l_um_iw[57] ;
 wire \top_I.branch[16].l_um_iw[58] ;
 wire \top_I.branch[16].l_um_iw[59] ;
 wire \top_I.branch[16].l_um_iw[5] ;
 wire \top_I.branch[16].l_um_iw[60] ;
 wire \top_I.branch[16].l_um_iw[61] ;
 wire \top_I.branch[16].l_um_iw[62] ;
 wire \top_I.branch[16].l_um_iw[63] ;
 wire \top_I.branch[16].l_um_iw[64] ;
 wire \top_I.branch[16].l_um_iw[65] ;
 wire \top_I.branch[16].l_um_iw[66] ;
 wire \top_I.branch[16].l_um_iw[67] ;
 wire \top_I.branch[16].l_um_iw[68] ;
 wire \top_I.branch[16].l_um_iw[69] ;
 wire \top_I.branch[16].l_um_iw[6] ;
 wire \top_I.branch[16].l_um_iw[70] ;
 wire \top_I.branch[16].l_um_iw[71] ;
 wire \top_I.branch[16].l_um_iw[72] ;
 wire \top_I.branch[16].l_um_iw[73] ;
 wire \top_I.branch[16].l_um_iw[74] ;
 wire \top_I.branch[16].l_um_iw[75] ;
 wire \top_I.branch[16].l_um_iw[76] ;
 wire \top_I.branch[16].l_um_iw[77] ;
 wire \top_I.branch[16].l_um_iw[78] ;
 wire \top_I.branch[16].l_um_iw[79] ;
 wire \top_I.branch[16].l_um_iw[7] ;
 wire \top_I.branch[16].l_um_iw[80] ;
 wire \top_I.branch[16].l_um_iw[81] ;
 wire \top_I.branch[16].l_um_iw[82] ;
 wire \top_I.branch[16].l_um_iw[83] ;
 wire \top_I.branch[16].l_um_iw[84] ;
 wire \top_I.branch[16].l_um_iw[85] ;
 wire \top_I.branch[16].l_um_iw[86] ;
 wire \top_I.branch[16].l_um_iw[87] ;
 wire \top_I.branch[16].l_um_iw[88] ;
 wire \top_I.branch[16].l_um_iw[89] ;
 wire \top_I.branch[16].l_um_iw[8] ;
 wire \top_I.branch[16].l_um_iw[90] ;
 wire \top_I.branch[16].l_um_iw[91] ;
 wire \top_I.branch[16].l_um_iw[92] ;
 wire \top_I.branch[16].l_um_iw[93] ;
 wire \top_I.branch[16].l_um_iw[94] ;
 wire \top_I.branch[16].l_um_iw[95] ;
 wire \top_I.branch[16].l_um_iw[96] ;
 wire \top_I.branch[16].l_um_iw[97] ;
 wire \top_I.branch[16].l_um_iw[98] ;
 wire \top_I.branch[16].l_um_iw[99] ;
 wire \top_I.branch[16].l_um_iw[9] ;
 wire \top_I.branch[16].l_um_k_zero[0] ;
 wire \top_I.branch[16].l_um_k_zero[10] ;
 wire \top_I.branch[16].l_um_k_zero[11] ;
 wire \top_I.branch[16].l_um_k_zero[12] ;
 wire \top_I.branch[16].l_um_k_zero[13] ;
 wire \top_I.branch[16].l_um_k_zero[14] ;
 wire \top_I.branch[16].l_um_k_zero[15] ;
 wire \top_I.branch[16].l_um_k_zero[1] ;
 wire \top_I.branch[16].l_um_k_zero[2] ;
 wire \top_I.branch[16].l_um_k_zero[3] ;
 wire \top_I.branch[16].l_um_k_zero[4] ;
 wire \top_I.branch[16].l_um_k_zero[5] ;
 wire \top_I.branch[16].l_um_k_zero[6] ;
 wire \top_I.branch[16].l_um_k_zero[7] ;
 wire \top_I.branch[16].l_um_k_zero[8] ;
 wire \top_I.branch[16].l_um_k_zero[9] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[17].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[17].l_k_one ;
 wire \top_I.branch[17].l_k_zero ;
 wire \top_I.branch[17].l_um_ena[0] ;
 wire \top_I.branch[17].l_um_ena[10] ;
 wire \top_I.branch[17].l_um_ena[11] ;
 wire \top_I.branch[17].l_um_ena[12] ;
 wire \top_I.branch[17].l_um_ena[13] ;
 wire \top_I.branch[17].l_um_ena[14] ;
 wire \top_I.branch[17].l_um_ena[15] ;
 wire \top_I.branch[17].l_um_ena[1] ;
 wire \top_I.branch[17].l_um_ena[2] ;
 wire \top_I.branch[17].l_um_ena[3] ;
 wire \top_I.branch[17].l_um_ena[4] ;
 wire \top_I.branch[17].l_um_ena[5] ;
 wire \top_I.branch[17].l_um_ena[6] ;
 wire \top_I.branch[17].l_um_ena[7] ;
 wire \top_I.branch[17].l_um_ena[8] ;
 wire \top_I.branch[17].l_um_ena[9] ;
 wire \top_I.branch[17].l_um_iw[0] ;
 wire \top_I.branch[17].l_um_iw[100] ;
 wire \top_I.branch[17].l_um_iw[101] ;
 wire \top_I.branch[17].l_um_iw[102] ;
 wire \top_I.branch[17].l_um_iw[103] ;
 wire \top_I.branch[17].l_um_iw[104] ;
 wire \top_I.branch[17].l_um_iw[105] ;
 wire \top_I.branch[17].l_um_iw[106] ;
 wire \top_I.branch[17].l_um_iw[107] ;
 wire \top_I.branch[17].l_um_iw[108] ;
 wire \top_I.branch[17].l_um_iw[109] ;
 wire \top_I.branch[17].l_um_iw[10] ;
 wire \top_I.branch[17].l_um_iw[110] ;
 wire \top_I.branch[17].l_um_iw[111] ;
 wire \top_I.branch[17].l_um_iw[112] ;
 wire \top_I.branch[17].l_um_iw[113] ;
 wire \top_I.branch[17].l_um_iw[114] ;
 wire \top_I.branch[17].l_um_iw[115] ;
 wire \top_I.branch[17].l_um_iw[116] ;
 wire \top_I.branch[17].l_um_iw[117] ;
 wire \top_I.branch[17].l_um_iw[118] ;
 wire \top_I.branch[17].l_um_iw[119] ;
 wire \top_I.branch[17].l_um_iw[11] ;
 wire \top_I.branch[17].l_um_iw[120] ;
 wire \top_I.branch[17].l_um_iw[121] ;
 wire \top_I.branch[17].l_um_iw[122] ;
 wire \top_I.branch[17].l_um_iw[123] ;
 wire \top_I.branch[17].l_um_iw[124] ;
 wire \top_I.branch[17].l_um_iw[125] ;
 wire \top_I.branch[17].l_um_iw[126] ;
 wire \top_I.branch[17].l_um_iw[127] ;
 wire \top_I.branch[17].l_um_iw[128] ;
 wire \top_I.branch[17].l_um_iw[129] ;
 wire \top_I.branch[17].l_um_iw[12] ;
 wire \top_I.branch[17].l_um_iw[130] ;
 wire \top_I.branch[17].l_um_iw[131] ;
 wire \top_I.branch[17].l_um_iw[132] ;
 wire \top_I.branch[17].l_um_iw[133] ;
 wire \top_I.branch[17].l_um_iw[134] ;
 wire \top_I.branch[17].l_um_iw[135] ;
 wire \top_I.branch[17].l_um_iw[136] ;
 wire \top_I.branch[17].l_um_iw[137] ;
 wire \top_I.branch[17].l_um_iw[138] ;
 wire \top_I.branch[17].l_um_iw[139] ;
 wire \top_I.branch[17].l_um_iw[13] ;
 wire \top_I.branch[17].l_um_iw[140] ;
 wire \top_I.branch[17].l_um_iw[141] ;
 wire \top_I.branch[17].l_um_iw[142] ;
 wire \top_I.branch[17].l_um_iw[143] ;
 wire \top_I.branch[17].l_um_iw[144] ;
 wire \top_I.branch[17].l_um_iw[145] ;
 wire \top_I.branch[17].l_um_iw[146] ;
 wire \top_I.branch[17].l_um_iw[147] ;
 wire \top_I.branch[17].l_um_iw[148] ;
 wire \top_I.branch[17].l_um_iw[149] ;
 wire \top_I.branch[17].l_um_iw[14] ;
 wire \top_I.branch[17].l_um_iw[150] ;
 wire \top_I.branch[17].l_um_iw[151] ;
 wire \top_I.branch[17].l_um_iw[152] ;
 wire \top_I.branch[17].l_um_iw[153] ;
 wire \top_I.branch[17].l_um_iw[154] ;
 wire \top_I.branch[17].l_um_iw[155] ;
 wire \top_I.branch[17].l_um_iw[156] ;
 wire \top_I.branch[17].l_um_iw[157] ;
 wire \top_I.branch[17].l_um_iw[158] ;
 wire \top_I.branch[17].l_um_iw[159] ;
 wire \top_I.branch[17].l_um_iw[15] ;
 wire \top_I.branch[17].l_um_iw[160] ;
 wire \top_I.branch[17].l_um_iw[161] ;
 wire \top_I.branch[17].l_um_iw[162] ;
 wire \top_I.branch[17].l_um_iw[163] ;
 wire \top_I.branch[17].l_um_iw[164] ;
 wire \top_I.branch[17].l_um_iw[165] ;
 wire \top_I.branch[17].l_um_iw[166] ;
 wire \top_I.branch[17].l_um_iw[167] ;
 wire \top_I.branch[17].l_um_iw[168] ;
 wire \top_I.branch[17].l_um_iw[169] ;
 wire \top_I.branch[17].l_um_iw[16] ;
 wire \top_I.branch[17].l_um_iw[170] ;
 wire \top_I.branch[17].l_um_iw[171] ;
 wire \top_I.branch[17].l_um_iw[172] ;
 wire \top_I.branch[17].l_um_iw[173] ;
 wire \top_I.branch[17].l_um_iw[174] ;
 wire \top_I.branch[17].l_um_iw[175] ;
 wire \top_I.branch[17].l_um_iw[176] ;
 wire \top_I.branch[17].l_um_iw[177] ;
 wire \top_I.branch[17].l_um_iw[178] ;
 wire \top_I.branch[17].l_um_iw[179] ;
 wire \top_I.branch[17].l_um_iw[17] ;
 wire \top_I.branch[17].l_um_iw[180] ;
 wire \top_I.branch[17].l_um_iw[181] ;
 wire \top_I.branch[17].l_um_iw[182] ;
 wire \top_I.branch[17].l_um_iw[183] ;
 wire \top_I.branch[17].l_um_iw[184] ;
 wire \top_I.branch[17].l_um_iw[185] ;
 wire \top_I.branch[17].l_um_iw[186] ;
 wire \top_I.branch[17].l_um_iw[187] ;
 wire \top_I.branch[17].l_um_iw[188] ;
 wire \top_I.branch[17].l_um_iw[189] ;
 wire \top_I.branch[17].l_um_iw[18] ;
 wire \top_I.branch[17].l_um_iw[190] ;
 wire \top_I.branch[17].l_um_iw[191] ;
 wire \top_I.branch[17].l_um_iw[192] ;
 wire \top_I.branch[17].l_um_iw[193] ;
 wire \top_I.branch[17].l_um_iw[194] ;
 wire \top_I.branch[17].l_um_iw[195] ;
 wire \top_I.branch[17].l_um_iw[196] ;
 wire \top_I.branch[17].l_um_iw[197] ;
 wire \top_I.branch[17].l_um_iw[198] ;
 wire \top_I.branch[17].l_um_iw[199] ;
 wire \top_I.branch[17].l_um_iw[19] ;
 wire \top_I.branch[17].l_um_iw[1] ;
 wire \top_I.branch[17].l_um_iw[200] ;
 wire \top_I.branch[17].l_um_iw[201] ;
 wire \top_I.branch[17].l_um_iw[202] ;
 wire \top_I.branch[17].l_um_iw[203] ;
 wire \top_I.branch[17].l_um_iw[204] ;
 wire \top_I.branch[17].l_um_iw[205] ;
 wire \top_I.branch[17].l_um_iw[206] ;
 wire \top_I.branch[17].l_um_iw[207] ;
 wire \top_I.branch[17].l_um_iw[208] ;
 wire \top_I.branch[17].l_um_iw[209] ;
 wire \top_I.branch[17].l_um_iw[20] ;
 wire \top_I.branch[17].l_um_iw[210] ;
 wire \top_I.branch[17].l_um_iw[211] ;
 wire \top_I.branch[17].l_um_iw[212] ;
 wire \top_I.branch[17].l_um_iw[213] ;
 wire \top_I.branch[17].l_um_iw[214] ;
 wire \top_I.branch[17].l_um_iw[215] ;
 wire \top_I.branch[17].l_um_iw[216] ;
 wire \top_I.branch[17].l_um_iw[217] ;
 wire \top_I.branch[17].l_um_iw[218] ;
 wire \top_I.branch[17].l_um_iw[219] ;
 wire \top_I.branch[17].l_um_iw[21] ;
 wire \top_I.branch[17].l_um_iw[220] ;
 wire \top_I.branch[17].l_um_iw[221] ;
 wire \top_I.branch[17].l_um_iw[222] ;
 wire \top_I.branch[17].l_um_iw[223] ;
 wire \top_I.branch[17].l_um_iw[224] ;
 wire \top_I.branch[17].l_um_iw[225] ;
 wire \top_I.branch[17].l_um_iw[226] ;
 wire \top_I.branch[17].l_um_iw[227] ;
 wire \top_I.branch[17].l_um_iw[228] ;
 wire \top_I.branch[17].l_um_iw[229] ;
 wire \top_I.branch[17].l_um_iw[22] ;
 wire \top_I.branch[17].l_um_iw[230] ;
 wire \top_I.branch[17].l_um_iw[231] ;
 wire \top_I.branch[17].l_um_iw[232] ;
 wire \top_I.branch[17].l_um_iw[233] ;
 wire \top_I.branch[17].l_um_iw[234] ;
 wire \top_I.branch[17].l_um_iw[235] ;
 wire \top_I.branch[17].l_um_iw[236] ;
 wire \top_I.branch[17].l_um_iw[237] ;
 wire \top_I.branch[17].l_um_iw[238] ;
 wire \top_I.branch[17].l_um_iw[239] ;
 wire \top_I.branch[17].l_um_iw[23] ;
 wire \top_I.branch[17].l_um_iw[240] ;
 wire \top_I.branch[17].l_um_iw[241] ;
 wire \top_I.branch[17].l_um_iw[242] ;
 wire \top_I.branch[17].l_um_iw[243] ;
 wire \top_I.branch[17].l_um_iw[244] ;
 wire \top_I.branch[17].l_um_iw[245] ;
 wire \top_I.branch[17].l_um_iw[246] ;
 wire \top_I.branch[17].l_um_iw[247] ;
 wire \top_I.branch[17].l_um_iw[248] ;
 wire \top_I.branch[17].l_um_iw[249] ;
 wire \top_I.branch[17].l_um_iw[24] ;
 wire \top_I.branch[17].l_um_iw[250] ;
 wire \top_I.branch[17].l_um_iw[251] ;
 wire \top_I.branch[17].l_um_iw[252] ;
 wire \top_I.branch[17].l_um_iw[253] ;
 wire \top_I.branch[17].l_um_iw[254] ;
 wire \top_I.branch[17].l_um_iw[255] ;
 wire \top_I.branch[17].l_um_iw[256] ;
 wire \top_I.branch[17].l_um_iw[257] ;
 wire \top_I.branch[17].l_um_iw[258] ;
 wire \top_I.branch[17].l_um_iw[259] ;
 wire \top_I.branch[17].l_um_iw[25] ;
 wire \top_I.branch[17].l_um_iw[260] ;
 wire \top_I.branch[17].l_um_iw[261] ;
 wire \top_I.branch[17].l_um_iw[262] ;
 wire \top_I.branch[17].l_um_iw[263] ;
 wire \top_I.branch[17].l_um_iw[264] ;
 wire \top_I.branch[17].l_um_iw[265] ;
 wire \top_I.branch[17].l_um_iw[266] ;
 wire \top_I.branch[17].l_um_iw[267] ;
 wire \top_I.branch[17].l_um_iw[268] ;
 wire \top_I.branch[17].l_um_iw[269] ;
 wire \top_I.branch[17].l_um_iw[26] ;
 wire \top_I.branch[17].l_um_iw[270] ;
 wire \top_I.branch[17].l_um_iw[271] ;
 wire \top_I.branch[17].l_um_iw[272] ;
 wire \top_I.branch[17].l_um_iw[273] ;
 wire \top_I.branch[17].l_um_iw[274] ;
 wire \top_I.branch[17].l_um_iw[275] ;
 wire \top_I.branch[17].l_um_iw[276] ;
 wire \top_I.branch[17].l_um_iw[277] ;
 wire \top_I.branch[17].l_um_iw[278] ;
 wire \top_I.branch[17].l_um_iw[279] ;
 wire \top_I.branch[17].l_um_iw[27] ;
 wire \top_I.branch[17].l_um_iw[280] ;
 wire \top_I.branch[17].l_um_iw[281] ;
 wire \top_I.branch[17].l_um_iw[282] ;
 wire \top_I.branch[17].l_um_iw[283] ;
 wire \top_I.branch[17].l_um_iw[284] ;
 wire \top_I.branch[17].l_um_iw[285] ;
 wire \top_I.branch[17].l_um_iw[286] ;
 wire \top_I.branch[17].l_um_iw[287] ;
 wire \top_I.branch[17].l_um_iw[28] ;
 wire \top_I.branch[17].l_um_iw[29] ;
 wire \top_I.branch[17].l_um_iw[2] ;
 wire \top_I.branch[17].l_um_iw[30] ;
 wire \top_I.branch[17].l_um_iw[31] ;
 wire \top_I.branch[17].l_um_iw[32] ;
 wire \top_I.branch[17].l_um_iw[33] ;
 wire \top_I.branch[17].l_um_iw[34] ;
 wire \top_I.branch[17].l_um_iw[35] ;
 wire \top_I.branch[17].l_um_iw[36] ;
 wire \top_I.branch[17].l_um_iw[37] ;
 wire \top_I.branch[17].l_um_iw[38] ;
 wire \top_I.branch[17].l_um_iw[39] ;
 wire \top_I.branch[17].l_um_iw[3] ;
 wire \top_I.branch[17].l_um_iw[40] ;
 wire \top_I.branch[17].l_um_iw[41] ;
 wire \top_I.branch[17].l_um_iw[42] ;
 wire \top_I.branch[17].l_um_iw[43] ;
 wire \top_I.branch[17].l_um_iw[44] ;
 wire \top_I.branch[17].l_um_iw[45] ;
 wire \top_I.branch[17].l_um_iw[46] ;
 wire \top_I.branch[17].l_um_iw[47] ;
 wire \top_I.branch[17].l_um_iw[48] ;
 wire \top_I.branch[17].l_um_iw[49] ;
 wire \top_I.branch[17].l_um_iw[4] ;
 wire \top_I.branch[17].l_um_iw[50] ;
 wire \top_I.branch[17].l_um_iw[51] ;
 wire \top_I.branch[17].l_um_iw[52] ;
 wire \top_I.branch[17].l_um_iw[53] ;
 wire \top_I.branch[17].l_um_iw[54] ;
 wire \top_I.branch[17].l_um_iw[55] ;
 wire \top_I.branch[17].l_um_iw[56] ;
 wire \top_I.branch[17].l_um_iw[57] ;
 wire \top_I.branch[17].l_um_iw[58] ;
 wire \top_I.branch[17].l_um_iw[59] ;
 wire \top_I.branch[17].l_um_iw[5] ;
 wire \top_I.branch[17].l_um_iw[60] ;
 wire \top_I.branch[17].l_um_iw[61] ;
 wire \top_I.branch[17].l_um_iw[62] ;
 wire \top_I.branch[17].l_um_iw[63] ;
 wire \top_I.branch[17].l_um_iw[64] ;
 wire \top_I.branch[17].l_um_iw[65] ;
 wire \top_I.branch[17].l_um_iw[66] ;
 wire \top_I.branch[17].l_um_iw[67] ;
 wire \top_I.branch[17].l_um_iw[68] ;
 wire \top_I.branch[17].l_um_iw[69] ;
 wire \top_I.branch[17].l_um_iw[6] ;
 wire \top_I.branch[17].l_um_iw[70] ;
 wire \top_I.branch[17].l_um_iw[71] ;
 wire \top_I.branch[17].l_um_iw[72] ;
 wire \top_I.branch[17].l_um_iw[73] ;
 wire \top_I.branch[17].l_um_iw[74] ;
 wire \top_I.branch[17].l_um_iw[75] ;
 wire \top_I.branch[17].l_um_iw[76] ;
 wire \top_I.branch[17].l_um_iw[77] ;
 wire \top_I.branch[17].l_um_iw[78] ;
 wire \top_I.branch[17].l_um_iw[79] ;
 wire \top_I.branch[17].l_um_iw[7] ;
 wire \top_I.branch[17].l_um_iw[80] ;
 wire \top_I.branch[17].l_um_iw[81] ;
 wire \top_I.branch[17].l_um_iw[82] ;
 wire \top_I.branch[17].l_um_iw[83] ;
 wire \top_I.branch[17].l_um_iw[84] ;
 wire \top_I.branch[17].l_um_iw[85] ;
 wire \top_I.branch[17].l_um_iw[86] ;
 wire \top_I.branch[17].l_um_iw[87] ;
 wire \top_I.branch[17].l_um_iw[88] ;
 wire \top_I.branch[17].l_um_iw[89] ;
 wire \top_I.branch[17].l_um_iw[8] ;
 wire \top_I.branch[17].l_um_iw[90] ;
 wire \top_I.branch[17].l_um_iw[91] ;
 wire \top_I.branch[17].l_um_iw[92] ;
 wire \top_I.branch[17].l_um_iw[93] ;
 wire \top_I.branch[17].l_um_iw[94] ;
 wire \top_I.branch[17].l_um_iw[95] ;
 wire \top_I.branch[17].l_um_iw[96] ;
 wire \top_I.branch[17].l_um_iw[97] ;
 wire \top_I.branch[17].l_um_iw[98] ;
 wire \top_I.branch[17].l_um_iw[99] ;
 wire \top_I.branch[17].l_um_iw[9] ;
 wire \top_I.branch[17].l_um_k_zero[0] ;
 wire \top_I.branch[17].l_um_k_zero[10] ;
 wire \top_I.branch[17].l_um_k_zero[11] ;
 wire \top_I.branch[17].l_um_k_zero[12] ;
 wire \top_I.branch[17].l_um_k_zero[13] ;
 wire \top_I.branch[17].l_um_k_zero[14] ;
 wire \top_I.branch[17].l_um_k_zero[15] ;
 wire \top_I.branch[17].l_um_k_zero[1] ;
 wire \top_I.branch[17].l_um_k_zero[2] ;
 wire \top_I.branch[17].l_um_k_zero[3] ;
 wire \top_I.branch[17].l_um_k_zero[4] ;
 wire \top_I.branch[17].l_um_k_zero[5] ;
 wire \top_I.branch[17].l_um_k_zero[6] ;
 wire \top_I.branch[17].l_um_k_zero[7] ;
 wire \top_I.branch[17].l_um_k_zero[8] ;
 wire \top_I.branch[17].l_um_k_zero[9] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[18].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[18].l_k_one ;
 wire \top_I.branch[18].l_k_zero ;
 wire \top_I.branch[18].l_um_ena[0] ;
 wire \top_I.branch[18].l_um_ena[10] ;
 wire \top_I.branch[18].l_um_ena[11] ;
 wire \top_I.branch[18].l_um_ena[12] ;
 wire \top_I.branch[18].l_um_ena[13] ;
 wire \top_I.branch[18].l_um_ena[14] ;
 wire \top_I.branch[18].l_um_ena[15] ;
 wire \top_I.branch[18].l_um_ena[1] ;
 wire \top_I.branch[18].l_um_ena[2] ;
 wire \top_I.branch[18].l_um_ena[3] ;
 wire \top_I.branch[18].l_um_ena[4] ;
 wire \top_I.branch[18].l_um_ena[5] ;
 wire \top_I.branch[18].l_um_ena[6] ;
 wire \top_I.branch[18].l_um_ena[7] ;
 wire \top_I.branch[18].l_um_ena[8] ;
 wire \top_I.branch[18].l_um_ena[9] ;
 wire \top_I.branch[18].l_um_iw[0] ;
 wire \top_I.branch[18].l_um_iw[100] ;
 wire \top_I.branch[18].l_um_iw[101] ;
 wire \top_I.branch[18].l_um_iw[102] ;
 wire \top_I.branch[18].l_um_iw[103] ;
 wire \top_I.branch[18].l_um_iw[104] ;
 wire \top_I.branch[18].l_um_iw[105] ;
 wire \top_I.branch[18].l_um_iw[106] ;
 wire \top_I.branch[18].l_um_iw[107] ;
 wire \top_I.branch[18].l_um_iw[108] ;
 wire \top_I.branch[18].l_um_iw[109] ;
 wire \top_I.branch[18].l_um_iw[10] ;
 wire \top_I.branch[18].l_um_iw[110] ;
 wire \top_I.branch[18].l_um_iw[111] ;
 wire \top_I.branch[18].l_um_iw[112] ;
 wire \top_I.branch[18].l_um_iw[113] ;
 wire \top_I.branch[18].l_um_iw[114] ;
 wire \top_I.branch[18].l_um_iw[115] ;
 wire \top_I.branch[18].l_um_iw[116] ;
 wire \top_I.branch[18].l_um_iw[117] ;
 wire \top_I.branch[18].l_um_iw[118] ;
 wire \top_I.branch[18].l_um_iw[119] ;
 wire \top_I.branch[18].l_um_iw[11] ;
 wire \top_I.branch[18].l_um_iw[120] ;
 wire \top_I.branch[18].l_um_iw[121] ;
 wire \top_I.branch[18].l_um_iw[122] ;
 wire \top_I.branch[18].l_um_iw[123] ;
 wire \top_I.branch[18].l_um_iw[124] ;
 wire \top_I.branch[18].l_um_iw[125] ;
 wire \top_I.branch[18].l_um_iw[126] ;
 wire \top_I.branch[18].l_um_iw[127] ;
 wire \top_I.branch[18].l_um_iw[128] ;
 wire \top_I.branch[18].l_um_iw[129] ;
 wire \top_I.branch[18].l_um_iw[12] ;
 wire \top_I.branch[18].l_um_iw[130] ;
 wire \top_I.branch[18].l_um_iw[131] ;
 wire \top_I.branch[18].l_um_iw[132] ;
 wire \top_I.branch[18].l_um_iw[133] ;
 wire \top_I.branch[18].l_um_iw[134] ;
 wire \top_I.branch[18].l_um_iw[135] ;
 wire \top_I.branch[18].l_um_iw[136] ;
 wire \top_I.branch[18].l_um_iw[137] ;
 wire \top_I.branch[18].l_um_iw[138] ;
 wire \top_I.branch[18].l_um_iw[139] ;
 wire \top_I.branch[18].l_um_iw[13] ;
 wire \top_I.branch[18].l_um_iw[140] ;
 wire \top_I.branch[18].l_um_iw[141] ;
 wire \top_I.branch[18].l_um_iw[142] ;
 wire \top_I.branch[18].l_um_iw[143] ;
 wire \top_I.branch[18].l_um_iw[144] ;
 wire \top_I.branch[18].l_um_iw[145] ;
 wire \top_I.branch[18].l_um_iw[146] ;
 wire \top_I.branch[18].l_um_iw[147] ;
 wire \top_I.branch[18].l_um_iw[148] ;
 wire \top_I.branch[18].l_um_iw[149] ;
 wire \top_I.branch[18].l_um_iw[14] ;
 wire \top_I.branch[18].l_um_iw[150] ;
 wire \top_I.branch[18].l_um_iw[151] ;
 wire \top_I.branch[18].l_um_iw[152] ;
 wire \top_I.branch[18].l_um_iw[153] ;
 wire \top_I.branch[18].l_um_iw[154] ;
 wire \top_I.branch[18].l_um_iw[155] ;
 wire \top_I.branch[18].l_um_iw[156] ;
 wire \top_I.branch[18].l_um_iw[157] ;
 wire \top_I.branch[18].l_um_iw[158] ;
 wire \top_I.branch[18].l_um_iw[159] ;
 wire \top_I.branch[18].l_um_iw[15] ;
 wire \top_I.branch[18].l_um_iw[160] ;
 wire \top_I.branch[18].l_um_iw[161] ;
 wire \top_I.branch[18].l_um_iw[162] ;
 wire \top_I.branch[18].l_um_iw[163] ;
 wire \top_I.branch[18].l_um_iw[164] ;
 wire \top_I.branch[18].l_um_iw[165] ;
 wire \top_I.branch[18].l_um_iw[166] ;
 wire \top_I.branch[18].l_um_iw[167] ;
 wire \top_I.branch[18].l_um_iw[168] ;
 wire \top_I.branch[18].l_um_iw[169] ;
 wire \top_I.branch[18].l_um_iw[16] ;
 wire \top_I.branch[18].l_um_iw[170] ;
 wire \top_I.branch[18].l_um_iw[171] ;
 wire \top_I.branch[18].l_um_iw[172] ;
 wire \top_I.branch[18].l_um_iw[173] ;
 wire \top_I.branch[18].l_um_iw[174] ;
 wire \top_I.branch[18].l_um_iw[175] ;
 wire \top_I.branch[18].l_um_iw[176] ;
 wire \top_I.branch[18].l_um_iw[177] ;
 wire \top_I.branch[18].l_um_iw[178] ;
 wire \top_I.branch[18].l_um_iw[179] ;
 wire \top_I.branch[18].l_um_iw[17] ;
 wire \top_I.branch[18].l_um_iw[180] ;
 wire \top_I.branch[18].l_um_iw[181] ;
 wire \top_I.branch[18].l_um_iw[182] ;
 wire \top_I.branch[18].l_um_iw[183] ;
 wire \top_I.branch[18].l_um_iw[184] ;
 wire \top_I.branch[18].l_um_iw[185] ;
 wire \top_I.branch[18].l_um_iw[186] ;
 wire \top_I.branch[18].l_um_iw[187] ;
 wire \top_I.branch[18].l_um_iw[188] ;
 wire \top_I.branch[18].l_um_iw[189] ;
 wire \top_I.branch[18].l_um_iw[18] ;
 wire \top_I.branch[18].l_um_iw[190] ;
 wire \top_I.branch[18].l_um_iw[191] ;
 wire \top_I.branch[18].l_um_iw[192] ;
 wire \top_I.branch[18].l_um_iw[193] ;
 wire \top_I.branch[18].l_um_iw[194] ;
 wire \top_I.branch[18].l_um_iw[195] ;
 wire \top_I.branch[18].l_um_iw[196] ;
 wire \top_I.branch[18].l_um_iw[197] ;
 wire \top_I.branch[18].l_um_iw[198] ;
 wire \top_I.branch[18].l_um_iw[199] ;
 wire \top_I.branch[18].l_um_iw[19] ;
 wire \top_I.branch[18].l_um_iw[1] ;
 wire \top_I.branch[18].l_um_iw[200] ;
 wire \top_I.branch[18].l_um_iw[201] ;
 wire \top_I.branch[18].l_um_iw[202] ;
 wire \top_I.branch[18].l_um_iw[203] ;
 wire \top_I.branch[18].l_um_iw[204] ;
 wire \top_I.branch[18].l_um_iw[205] ;
 wire \top_I.branch[18].l_um_iw[206] ;
 wire \top_I.branch[18].l_um_iw[207] ;
 wire \top_I.branch[18].l_um_iw[208] ;
 wire \top_I.branch[18].l_um_iw[209] ;
 wire \top_I.branch[18].l_um_iw[20] ;
 wire \top_I.branch[18].l_um_iw[210] ;
 wire \top_I.branch[18].l_um_iw[211] ;
 wire \top_I.branch[18].l_um_iw[212] ;
 wire \top_I.branch[18].l_um_iw[213] ;
 wire \top_I.branch[18].l_um_iw[214] ;
 wire \top_I.branch[18].l_um_iw[215] ;
 wire \top_I.branch[18].l_um_iw[216] ;
 wire \top_I.branch[18].l_um_iw[217] ;
 wire \top_I.branch[18].l_um_iw[218] ;
 wire \top_I.branch[18].l_um_iw[219] ;
 wire \top_I.branch[18].l_um_iw[21] ;
 wire \top_I.branch[18].l_um_iw[220] ;
 wire \top_I.branch[18].l_um_iw[221] ;
 wire \top_I.branch[18].l_um_iw[222] ;
 wire \top_I.branch[18].l_um_iw[223] ;
 wire \top_I.branch[18].l_um_iw[224] ;
 wire \top_I.branch[18].l_um_iw[225] ;
 wire \top_I.branch[18].l_um_iw[226] ;
 wire \top_I.branch[18].l_um_iw[227] ;
 wire \top_I.branch[18].l_um_iw[228] ;
 wire \top_I.branch[18].l_um_iw[229] ;
 wire \top_I.branch[18].l_um_iw[22] ;
 wire \top_I.branch[18].l_um_iw[230] ;
 wire \top_I.branch[18].l_um_iw[231] ;
 wire \top_I.branch[18].l_um_iw[232] ;
 wire \top_I.branch[18].l_um_iw[233] ;
 wire \top_I.branch[18].l_um_iw[234] ;
 wire \top_I.branch[18].l_um_iw[235] ;
 wire \top_I.branch[18].l_um_iw[236] ;
 wire \top_I.branch[18].l_um_iw[237] ;
 wire \top_I.branch[18].l_um_iw[238] ;
 wire \top_I.branch[18].l_um_iw[239] ;
 wire \top_I.branch[18].l_um_iw[23] ;
 wire \top_I.branch[18].l_um_iw[240] ;
 wire \top_I.branch[18].l_um_iw[241] ;
 wire \top_I.branch[18].l_um_iw[242] ;
 wire \top_I.branch[18].l_um_iw[243] ;
 wire \top_I.branch[18].l_um_iw[244] ;
 wire \top_I.branch[18].l_um_iw[245] ;
 wire \top_I.branch[18].l_um_iw[246] ;
 wire \top_I.branch[18].l_um_iw[247] ;
 wire \top_I.branch[18].l_um_iw[248] ;
 wire \top_I.branch[18].l_um_iw[249] ;
 wire \top_I.branch[18].l_um_iw[24] ;
 wire \top_I.branch[18].l_um_iw[250] ;
 wire \top_I.branch[18].l_um_iw[251] ;
 wire \top_I.branch[18].l_um_iw[252] ;
 wire \top_I.branch[18].l_um_iw[253] ;
 wire \top_I.branch[18].l_um_iw[254] ;
 wire \top_I.branch[18].l_um_iw[255] ;
 wire \top_I.branch[18].l_um_iw[256] ;
 wire \top_I.branch[18].l_um_iw[257] ;
 wire \top_I.branch[18].l_um_iw[258] ;
 wire \top_I.branch[18].l_um_iw[259] ;
 wire \top_I.branch[18].l_um_iw[25] ;
 wire \top_I.branch[18].l_um_iw[260] ;
 wire \top_I.branch[18].l_um_iw[261] ;
 wire \top_I.branch[18].l_um_iw[262] ;
 wire \top_I.branch[18].l_um_iw[263] ;
 wire \top_I.branch[18].l_um_iw[264] ;
 wire \top_I.branch[18].l_um_iw[265] ;
 wire \top_I.branch[18].l_um_iw[266] ;
 wire \top_I.branch[18].l_um_iw[267] ;
 wire \top_I.branch[18].l_um_iw[268] ;
 wire \top_I.branch[18].l_um_iw[269] ;
 wire \top_I.branch[18].l_um_iw[26] ;
 wire \top_I.branch[18].l_um_iw[270] ;
 wire \top_I.branch[18].l_um_iw[271] ;
 wire \top_I.branch[18].l_um_iw[272] ;
 wire \top_I.branch[18].l_um_iw[273] ;
 wire \top_I.branch[18].l_um_iw[274] ;
 wire \top_I.branch[18].l_um_iw[275] ;
 wire \top_I.branch[18].l_um_iw[276] ;
 wire \top_I.branch[18].l_um_iw[277] ;
 wire \top_I.branch[18].l_um_iw[278] ;
 wire \top_I.branch[18].l_um_iw[279] ;
 wire \top_I.branch[18].l_um_iw[27] ;
 wire \top_I.branch[18].l_um_iw[280] ;
 wire \top_I.branch[18].l_um_iw[281] ;
 wire \top_I.branch[18].l_um_iw[282] ;
 wire \top_I.branch[18].l_um_iw[283] ;
 wire \top_I.branch[18].l_um_iw[284] ;
 wire \top_I.branch[18].l_um_iw[285] ;
 wire \top_I.branch[18].l_um_iw[286] ;
 wire \top_I.branch[18].l_um_iw[287] ;
 wire \top_I.branch[18].l_um_iw[28] ;
 wire \top_I.branch[18].l_um_iw[29] ;
 wire \top_I.branch[18].l_um_iw[2] ;
 wire \top_I.branch[18].l_um_iw[30] ;
 wire \top_I.branch[18].l_um_iw[31] ;
 wire \top_I.branch[18].l_um_iw[32] ;
 wire \top_I.branch[18].l_um_iw[33] ;
 wire \top_I.branch[18].l_um_iw[34] ;
 wire \top_I.branch[18].l_um_iw[35] ;
 wire \top_I.branch[18].l_um_iw[36] ;
 wire \top_I.branch[18].l_um_iw[37] ;
 wire \top_I.branch[18].l_um_iw[38] ;
 wire \top_I.branch[18].l_um_iw[39] ;
 wire \top_I.branch[18].l_um_iw[3] ;
 wire \top_I.branch[18].l_um_iw[40] ;
 wire \top_I.branch[18].l_um_iw[41] ;
 wire \top_I.branch[18].l_um_iw[42] ;
 wire \top_I.branch[18].l_um_iw[43] ;
 wire \top_I.branch[18].l_um_iw[44] ;
 wire \top_I.branch[18].l_um_iw[45] ;
 wire \top_I.branch[18].l_um_iw[46] ;
 wire \top_I.branch[18].l_um_iw[47] ;
 wire \top_I.branch[18].l_um_iw[48] ;
 wire \top_I.branch[18].l_um_iw[49] ;
 wire \top_I.branch[18].l_um_iw[4] ;
 wire \top_I.branch[18].l_um_iw[50] ;
 wire \top_I.branch[18].l_um_iw[51] ;
 wire \top_I.branch[18].l_um_iw[52] ;
 wire \top_I.branch[18].l_um_iw[53] ;
 wire \top_I.branch[18].l_um_iw[54] ;
 wire \top_I.branch[18].l_um_iw[55] ;
 wire \top_I.branch[18].l_um_iw[56] ;
 wire \top_I.branch[18].l_um_iw[57] ;
 wire \top_I.branch[18].l_um_iw[58] ;
 wire \top_I.branch[18].l_um_iw[59] ;
 wire \top_I.branch[18].l_um_iw[5] ;
 wire \top_I.branch[18].l_um_iw[60] ;
 wire \top_I.branch[18].l_um_iw[61] ;
 wire \top_I.branch[18].l_um_iw[62] ;
 wire \top_I.branch[18].l_um_iw[63] ;
 wire \top_I.branch[18].l_um_iw[64] ;
 wire \top_I.branch[18].l_um_iw[65] ;
 wire \top_I.branch[18].l_um_iw[66] ;
 wire \top_I.branch[18].l_um_iw[67] ;
 wire \top_I.branch[18].l_um_iw[68] ;
 wire \top_I.branch[18].l_um_iw[69] ;
 wire \top_I.branch[18].l_um_iw[6] ;
 wire \top_I.branch[18].l_um_iw[70] ;
 wire \top_I.branch[18].l_um_iw[71] ;
 wire \top_I.branch[18].l_um_iw[72] ;
 wire \top_I.branch[18].l_um_iw[73] ;
 wire \top_I.branch[18].l_um_iw[74] ;
 wire \top_I.branch[18].l_um_iw[75] ;
 wire \top_I.branch[18].l_um_iw[76] ;
 wire \top_I.branch[18].l_um_iw[77] ;
 wire \top_I.branch[18].l_um_iw[78] ;
 wire \top_I.branch[18].l_um_iw[79] ;
 wire \top_I.branch[18].l_um_iw[7] ;
 wire \top_I.branch[18].l_um_iw[80] ;
 wire \top_I.branch[18].l_um_iw[81] ;
 wire \top_I.branch[18].l_um_iw[82] ;
 wire \top_I.branch[18].l_um_iw[83] ;
 wire \top_I.branch[18].l_um_iw[84] ;
 wire \top_I.branch[18].l_um_iw[85] ;
 wire \top_I.branch[18].l_um_iw[86] ;
 wire \top_I.branch[18].l_um_iw[87] ;
 wire \top_I.branch[18].l_um_iw[88] ;
 wire \top_I.branch[18].l_um_iw[89] ;
 wire \top_I.branch[18].l_um_iw[8] ;
 wire \top_I.branch[18].l_um_iw[90] ;
 wire \top_I.branch[18].l_um_iw[91] ;
 wire \top_I.branch[18].l_um_iw[92] ;
 wire \top_I.branch[18].l_um_iw[93] ;
 wire \top_I.branch[18].l_um_iw[94] ;
 wire \top_I.branch[18].l_um_iw[95] ;
 wire \top_I.branch[18].l_um_iw[96] ;
 wire \top_I.branch[18].l_um_iw[97] ;
 wire \top_I.branch[18].l_um_iw[98] ;
 wire \top_I.branch[18].l_um_iw[99] ;
 wire \top_I.branch[18].l_um_iw[9] ;
 wire \top_I.branch[18].l_um_k_zero[0] ;
 wire \top_I.branch[18].l_um_k_zero[10] ;
 wire \top_I.branch[18].l_um_k_zero[11] ;
 wire \top_I.branch[18].l_um_k_zero[12] ;
 wire \top_I.branch[18].l_um_k_zero[13] ;
 wire \top_I.branch[18].l_um_k_zero[14] ;
 wire \top_I.branch[18].l_um_k_zero[15] ;
 wire \top_I.branch[18].l_um_k_zero[1] ;
 wire \top_I.branch[18].l_um_k_zero[2] ;
 wire \top_I.branch[18].l_um_k_zero[3] ;
 wire \top_I.branch[18].l_um_k_zero[4] ;
 wire \top_I.branch[18].l_um_k_zero[5] ;
 wire \top_I.branch[18].l_um_k_zero[6] ;
 wire \top_I.branch[18].l_um_k_zero[7] ;
 wire \top_I.branch[18].l_um_k_zero[8] ;
 wire \top_I.branch[18].l_um_k_zero[9] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[19].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[19].l_k_one ;
 wire \top_I.branch[19].l_k_zero ;
 wire \top_I.branch[19].l_um_ena[0] ;
 wire \top_I.branch[19].l_um_ena[10] ;
 wire \top_I.branch[19].l_um_ena[11] ;
 wire \top_I.branch[19].l_um_ena[12] ;
 wire \top_I.branch[19].l_um_ena[13] ;
 wire \top_I.branch[19].l_um_ena[14] ;
 wire \top_I.branch[19].l_um_ena[15] ;
 wire \top_I.branch[19].l_um_ena[1] ;
 wire \top_I.branch[19].l_um_ena[2] ;
 wire \top_I.branch[19].l_um_ena[3] ;
 wire \top_I.branch[19].l_um_ena[4] ;
 wire \top_I.branch[19].l_um_ena[5] ;
 wire \top_I.branch[19].l_um_ena[6] ;
 wire \top_I.branch[19].l_um_ena[7] ;
 wire \top_I.branch[19].l_um_ena[8] ;
 wire \top_I.branch[19].l_um_ena[9] ;
 wire \top_I.branch[19].l_um_iw[0] ;
 wire \top_I.branch[19].l_um_iw[100] ;
 wire \top_I.branch[19].l_um_iw[101] ;
 wire \top_I.branch[19].l_um_iw[102] ;
 wire \top_I.branch[19].l_um_iw[103] ;
 wire \top_I.branch[19].l_um_iw[104] ;
 wire \top_I.branch[19].l_um_iw[105] ;
 wire \top_I.branch[19].l_um_iw[106] ;
 wire \top_I.branch[19].l_um_iw[107] ;
 wire \top_I.branch[19].l_um_iw[108] ;
 wire \top_I.branch[19].l_um_iw[109] ;
 wire \top_I.branch[19].l_um_iw[10] ;
 wire \top_I.branch[19].l_um_iw[110] ;
 wire \top_I.branch[19].l_um_iw[111] ;
 wire \top_I.branch[19].l_um_iw[112] ;
 wire \top_I.branch[19].l_um_iw[113] ;
 wire \top_I.branch[19].l_um_iw[114] ;
 wire \top_I.branch[19].l_um_iw[115] ;
 wire \top_I.branch[19].l_um_iw[116] ;
 wire \top_I.branch[19].l_um_iw[117] ;
 wire \top_I.branch[19].l_um_iw[118] ;
 wire \top_I.branch[19].l_um_iw[119] ;
 wire \top_I.branch[19].l_um_iw[11] ;
 wire \top_I.branch[19].l_um_iw[120] ;
 wire \top_I.branch[19].l_um_iw[121] ;
 wire \top_I.branch[19].l_um_iw[122] ;
 wire \top_I.branch[19].l_um_iw[123] ;
 wire \top_I.branch[19].l_um_iw[124] ;
 wire \top_I.branch[19].l_um_iw[125] ;
 wire \top_I.branch[19].l_um_iw[126] ;
 wire \top_I.branch[19].l_um_iw[127] ;
 wire \top_I.branch[19].l_um_iw[128] ;
 wire \top_I.branch[19].l_um_iw[129] ;
 wire \top_I.branch[19].l_um_iw[12] ;
 wire \top_I.branch[19].l_um_iw[130] ;
 wire \top_I.branch[19].l_um_iw[131] ;
 wire \top_I.branch[19].l_um_iw[132] ;
 wire \top_I.branch[19].l_um_iw[133] ;
 wire \top_I.branch[19].l_um_iw[134] ;
 wire \top_I.branch[19].l_um_iw[135] ;
 wire \top_I.branch[19].l_um_iw[136] ;
 wire \top_I.branch[19].l_um_iw[137] ;
 wire \top_I.branch[19].l_um_iw[138] ;
 wire \top_I.branch[19].l_um_iw[139] ;
 wire \top_I.branch[19].l_um_iw[13] ;
 wire \top_I.branch[19].l_um_iw[140] ;
 wire \top_I.branch[19].l_um_iw[141] ;
 wire \top_I.branch[19].l_um_iw[142] ;
 wire \top_I.branch[19].l_um_iw[143] ;
 wire \top_I.branch[19].l_um_iw[144] ;
 wire \top_I.branch[19].l_um_iw[145] ;
 wire \top_I.branch[19].l_um_iw[146] ;
 wire \top_I.branch[19].l_um_iw[147] ;
 wire \top_I.branch[19].l_um_iw[148] ;
 wire \top_I.branch[19].l_um_iw[149] ;
 wire \top_I.branch[19].l_um_iw[14] ;
 wire \top_I.branch[19].l_um_iw[150] ;
 wire \top_I.branch[19].l_um_iw[151] ;
 wire \top_I.branch[19].l_um_iw[152] ;
 wire \top_I.branch[19].l_um_iw[153] ;
 wire \top_I.branch[19].l_um_iw[154] ;
 wire \top_I.branch[19].l_um_iw[155] ;
 wire \top_I.branch[19].l_um_iw[156] ;
 wire \top_I.branch[19].l_um_iw[157] ;
 wire \top_I.branch[19].l_um_iw[158] ;
 wire \top_I.branch[19].l_um_iw[159] ;
 wire \top_I.branch[19].l_um_iw[15] ;
 wire \top_I.branch[19].l_um_iw[160] ;
 wire \top_I.branch[19].l_um_iw[161] ;
 wire \top_I.branch[19].l_um_iw[162] ;
 wire \top_I.branch[19].l_um_iw[163] ;
 wire \top_I.branch[19].l_um_iw[164] ;
 wire \top_I.branch[19].l_um_iw[165] ;
 wire \top_I.branch[19].l_um_iw[166] ;
 wire \top_I.branch[19].l_um_iw[167] ;
 wire \top_I.branch[19].l_um_iw[168] ;
 wire \top_I.branch[19].l_um_iw[169] ;
 wire \top_I.branch[19].l_um_iw[16] ;
 wire \top_I.branch[19].l_um_iw[170] ;
 wire \top_I.branch[19].l_um_iw[171] ;
 wire \top_I.branch[19].l_um_iw[172] ;
 wire \top_I.branch[19].l_um_iw[173] ;
 wire \top_I.branch[19].l_um_iw[174] ;
 wire \top_I.branch[19].l_um_iw[175] ;
 wire \top_I.branch[19].l_um_iw[176] ;
 wire \top_I.branch[19].l_um_iw[177] ;
 wire \top_I.branch[19].l_um_iw[178] ;
 wire \top_I.branch[19].l_um_iw[179] ;
 wire \top_I.branch[19].l_um_iw[17] ;
 wire \top_I.branch[19].l_um_iw[180] ;
 wire \top_I.branch[19].l_um_iw[181] ;
 wire \top_I.branch[19].l_um_iw[182] ;
 wire \top_I.branch[19].l_um_iw[183] ;
 wire \top_I.branch[19].l_um_iw[184] ;
 wire \top_I.branch[19].l_um_iw[185] ;
 wire \top_I.branch[19].l_um_iw[186] ;
 wire \top_I.branch[19].l_um_iw[187] ;
 wire \top_I.branch[19].l_um_iw[188] ;
 wire \top_I.branch[19].l_um_iw[189] ;
 wire \top_I.branch[19].l_um_iw[18] ;
 wire \top_I.branch[19].l_um_iw[190] ;
 wire \top_I.branch[19].l_um_iw[191] ;
 wire \top_I.branch[19].l_um_iw[192] ;
 wire \top_I.branch[19].l_um_iw[193] ;
 wire \top_I.branch[19].l_um_iw[194] ;
 wire \top_I.branch[19].l_um_iw[195] ;
 wire \top_I.branch[19].l_um_iw[196] ;
 wire \top_I.branch[19].l_um_iw[197] ;
 wire \top_I.branch[19].l_um_iw[198] ;
 wire \top_I.branch[19].l_um_iw[199] ;
 wire \top_I.branch[19].l_um_iw[19] ;
 wire \top_I.branch[19].l_um_iw[1] ;
 wire \top_I.branch[19].l_um_iw[200] ;
 wire \top_I.branch[19].l_um_iw[201] ;
 wire \top_I.branch[19].l_um_iw[202] ;
 wire \top_I.branch[19].l_um_iw[203] ;
 wire \top_I.branch[19].l_um_iw[204] ;
 wire \top_I.branch[19].l_um_iw[205] ;
 wire \top_I.branch[19].l_um_iw[206] ;
 wire \top_I.branch[19].l_um_iw[207] ;
 wire \top_I.branch[19].l_um_iw[208] ;
 wire \top_I.branch[19].l_um_iw[209] ;
 wire \top_I.branch[19].l_um_iw[20] ;
 wire \top_I.branch[19].l_um_iw[210] ;
 wire \top_I.branch[19].l_um_iw[211] ;
 wire \top_I.branch[19].l_um_iw[212] ;
 wire \top_I.branch[19].l_um_iw[213] ;
 wire \top_I.branch[19].l_um_iw[214] ;
 wire \top_I.branch[19].l_um_iw[215] ;
 wire \top_I.branch[19].l_um_iw[216] ;
 wire \top_I.branch[19].l_um_iw[217] ;
 wire \top_I.branch[19].l_um_iw[218] ;
 wire \top_I.branch[19].l_um_iw[219] ;
 wire \top_I.branch[19].l_um_iw[21] ;
 wire \top_I.branch[19].l_um_iw[220] ;
 wire \top_I.branch[19].l_um_iw[221] ;
 wire \top_I.branch[19].l_um_iw[222] ;
 wire \top_I.branch[19].l_um_iw[223] ;
 wire \top_I.branch[19].l_um_iw[224] ;
 wire \top_I.branch[19].l_um_iw[225] ;
 wire \top_I.branch[19].l_um_iw[226] ;
 wire \top_I.branch[19].l_um_iw[227] ;
 wire \top_I.branch[19].l_um_iw[228] ;
 wire \top_I.branch[19].l_um_iw[229] ;
 wire \top_I.branch[19].l_um_iw[22] ;
 wire \top_I.branch[19].l_um_iw[230] ;
 wire \top_I.branch[19].l_um_iw[231] ;
 wire \top_I.branch[19].l_um_iw[232] ;
 wire \top_I.branch[19].l_um_iw[233] ;
 wire \top_I.branch[19].l_um_iw[234] ;
 wire \top_I.branch[19].l_um_iw[235] ;
 wire \top_I.branch[19].l_um_iw[236] ;
 wire \top_I.branch[19].l_um_iw[237] ;
 wire \top_I.branch[19].l_um_iw[238] ;
 wire \top_I.branch[19].l_um_iw[239] ;
 wire \top_I.branch[19].l_um_iw[23] ;
 wire \top_I.branch[19].l_um_iw[240] ;
 wire \top_I.branch[19].l_um_iw[241] ;
 wire \top_I.branch[19].l_um_iw[242] ;
 wire \top_I.branch[19].l_um_iw[243] ;
 wire \top_I.branch[19].l_um_iw[244] ;
 wire \top_I.branch[19].l_um_iw[245] ;
 wire \top_I.branch[19].l_um_iw[246] ;
 wire \top_I.branch[19].l_um_iw[247] ;
 wire \top_I.branch[19].l_um_iw[248] ;
 wire \top_I.branch[19].l_um_iw[249] ;
 wire \top_I.branch[19].l_um_iw[24] ;
 wire \top_I.branch[19].l_um_iw[250] ;
 wire \top_I.branch[19].l_um_iw[251] ;
 wire \top_I.branch[19].l_um_iw[252] ;
 wire \top_I.branch[19].l_um_iw[253] ;
 wire \top_I.branch[19].l_um_iw[254] ;
 wire \top_I.branch[19].l_um_iw[255] ;
 wire \top_I.branch[19].l_um_iw[256] ;
 wire \top_I.branch[19].l_um_iw[257] ;
 wire \top_I.branch[19].l_um_iw[258] ;
 wire \top_I.branch[19].l_um_iw[259] ;
 wire \top_I.branch[19].l_um_iw[25] ;
 wire \top_I.branch[19].l_um_iw[260] ;
 wire \top_I.branch[19].l_um_iw[261] ;
 wire \top_I.branch[19].l_um_iw[262] ;
 wire \top_I.branch[19].l_um_iw[263] ;
 wire \top_I.branch[19].l_um_iw[264] ;
 wire \top_I.branch[19].l_um_iw[265] ;
 wire \top_I.branch[19].l_um_iw[266] ;
 wire \top_I.branch[19].l_um_iw[267] ;
 wire \top_I.branch[19].l_um_iw[268] ;
 wire \top_I.branch[19].l_um_iw[269] ;
 wire \top_I.branch[19].l_um_iw[26] ;
 wire \top_I.branch[19].l_um_iw[270] ;
 wire \top_I.branch[19].l_um_iw[271] ;
 wire \top_I.branch[19].l_um_iw[272] ;
 wire \top_I.branch[19].l_um_iw[273] ;
 wire \top_I.branch[19].l_um_iw[274] ;
 wire \top_I.branch[19].l_um_iw[275] ;
 wire \top_I.branch[19].l_um_iw[276] ;
 wire \top_I.branch[19].l_um_iw[277] ;
 wire \top_I.branch[19].l_um_iw[278] ;
 wire \top_I.branch[19].l_um_iw[279] ;
 wire \top_I.branch[19].l_um_iw[27] ;
 wire \top_I.branch[19].l_um_iw[280] ;
 wire \top_I.branch[19].l_um_iw[281] ;
 wire \top_I.branch[19].l_um_iw[282] ;
 wire \top_I.branch[19].l_um_iw[283] ;
 wire \top_I.branch[19].l_um_iw[284] ;
 wire \top_I.branch[19].l_um_iw[285] ;
 wire \top_I.branch[19].l_um_iw[286] ;
 wire \top_I.branch[19].l_um_iw[287] ;
 wire \top_I.branch[19].l_um_iw[28] ;
 wire \top_I.branch[19].l_um_iw[29] ;
 wire \top_I.branch[19].l_um_iw[2] ;
 wire \top_I.branch[19].l_um_iw[30] ;
 wire \top_I.branch[19].l_um_iw[31] ;
 wire \top_I.branch[19].l_um_iw[32] ;
 wire \top_I.branch[19].l_um_iw[33] ;
 wire \top_I.branch[19].l_um_iw[34] ;
 wire \top_I.branch[19].l_um_iw[35] ;
 wire \top_I.branch[19].l_um_iw[36] ;
 wire \top_I.branch[19].l_um_iw[37] ;
 wire \top_I.branch[19].l_um_iw[38] ;
 wire \top_I.branch[19].l_um_iw[39] ;
 wire \top_I.branch[19].l_um_iw[3] ;
 wire \top_I.branch[19].l_um_iw[40] ;
 wire \top_I.branch[19].l_um_iw[41] ;
 wire \top_I.branch[19].l_um_iw[42] ;
 wire \top_I.branch[19].l_um_iw[43] ;
 wire \top_I.branch[19].l_um_iw[44] ;
 wire \top_I.branch[19].l_um_iw[45] ;
 wire \top_I.branch[19].l_um_iw[46] ;
 wire \top_I.branch[19].l_um_iw[47] ;
 wire \top_I.branch[19].l_um_iw[48] ;
 wire \top_I.branch[19].l_um_iw[49] ;
 wire \top_I.branch[19].l_um_iw[4] ;
 wire \top_I.branch[19].l_um_iw[50] ;
 wire \top_I.branch[19].l_um_iw[51] ;
 wire \top_I.branch[19].l_um_iw[52] ;
 wire \top_I.branch[19].l_um_iw[53] ;
 wire \top_I.branch[19].l_um_iw[54] ;
 wire \top_I.branch[19].l_um_iw[55] ;
 wire \top_I.branch[19].l_um_iw[56] ;
 wire \top_I.branch[19].l_um_iw[57] ;
 wire \top_I.branch[19].l_um_iw[58] ;
 wire \top_I.branch[19].l_um_iw[59] ;
 wire \top_I.branch[19].l_um_iw[5] ;
 wire \top_I.branch[19].l_um_iw[60] ;
 wire \top_I.branch[19].l_um_iw[61] ;
 wire \top_I.branch[19].l_um_iw[62] ;
 wire \top_I.branch[19].l_um_iw[63] ;
 wire \top_I.branch[19].l_um_iw[64] ;
 wire \top_I.branch[19].l_um_iw[65] ;
 wire \top_I.branch[19].l_um_iw[66] ;
 wire \top_I.branch[19].l_um_iw[67] ;
 wire \top_I.branch[19].l_um_iw[68] ;
 wire \top_I.branch[19].l_um_iw[69] ;
 wire \top_I.branch[19].l_um_iw[6] ;
 wire \top_I.branch[19].l_um_iw[70] ;
 wire \top_I.branch[19].l_um_iw[71] ;
 wire \top_I.branch[19].l_um_iw[72] ;
 wire \top_I.branch[19].l_um_iw[73] ;
 wire \top_I.branch[19].l_um_iw[74] ;
 wire \top_I.branch[19].l_um_iw[75] ;
 wire \top_I.branch[19].l_um_iw[76] ;
 wire \top_I.branch[19].l_um_iw[77] ;
 wire \top_I.branch[19].l_um_iw[78] ;
 wire \top_I.branch[19].l_um_iw[79] ;
 wire \top_I.branch[19].l_um_iw[7] ;
 wire \top_I.branch[19].l_um_iw[80] ;
 wire \top_I.branch[19].l_um_iw[81] ;
 wire \top_I.branch[19].l_um_iw[82] ;
 wire \top_I.branch[19].l_um_iw[83] ;
 wire \top_I.branch[19].l_um_iw[84] ;
 wire \top_I.branch[19].l_um_iw[85] ;
 wire \top_I.branch[19].l_um_iw[86] ;
 wire \top_I.branch[19].l_um_iw[87] ;
 wire \top_I.branch[19].l_um_iw[88] ;
 wire \top_I.branch[19].l_um_iw[89] ;
 wire \top_I.branch[19].l_um_iw[8] ;
 wire \top_I.branch[19].l_um_iw[90] ;
 wire \top_I.branch[19].l_um_iw[91] ;
 wire \top_I.branch[19].l_um_iw[92] ;
 wire \top_I.branch[19].l_um_iw[93] ;
 wire \top_I.branch[19].l_um_iw[94] ;
 wire \top_I.branch[19].l_um_iw[95] ;
 wire \top_I.branch[19].l_um_iw[96] ;
 wire \top_I.branch[19].l_um_iw[97] ;
 wire \top_I.branch[19].l_um_iw[98] ;
 wire \top_I.branch[19].l_um_iw[99] ;
 wire \top_I.branch[19].l_um_iw[9] ;
 wire \top_I.branch[19].l_um_k_zero[0] ;
 wire \top_I.branch[19].l_um_k_zero[10] ;
 wire \top_I.branch[19].l_um_k_zero[11] ;
 wire \top_I.branch[19].l_um_k_zero[12] ;
 wire \top_I.branch[19].l_um_k_zero[13] ;
 wire \top_I.branch[19].l_um_k_zero[14] ;
 wire \top_I.branch[19].l_um_k_zero[15] ;
 wire \top_I.branch[19].l_um_k_zero[1] ;
 wire \top_I.branch[19].l_um_k_zero[2] ;
 wire \top_I.branch[19].l_um_k_zero[3] ;
 wire \top_I.branch[19].l_um_k_zero[4] ;
 wire \top_I.branch[19].l_um_k_zero[5] ;
 wire \top_I.branch[19].l_um_k_zero[6] ;
 wire \top_I.branch[19].l_um_k_zero[7] ;
 wire \top_I.branch[19].l_um_k_zero[8] ;
 wire \top_I.branch[19].l_um_k_zero[9] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[1].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[2].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[2].um_top_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[3].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[4].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[4].um_top_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[5].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[6].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[6].um_top_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[7].um_bot_I.uo_out[7] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[0] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[1] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[2] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[3] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[4] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[5] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[6] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_oe[7] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[0] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[1] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[2] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[3] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[4] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[5] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[6] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uio_out[7] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[0] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[1] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[2] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[3] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[4] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[5] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[6] ;
 wire \top_I.branch[1].col_um[7].um_top_I.uo_out[7] ;
 wire \top_I.branch[1].l_k_one ;
 wire \top_I.branch[1].l_k_zero ;
 wire \top_I.branch[1].l_um_ena[0] ;
 wire \top_I.branch[1].l_um_ena[10] ;
 wire \top_I.branch[1].l_um_ena[11] ;
 wire \top_I.branch[1].l_um_ena[12] ;
 wire \top_I.branch[1].l_um_ena[13] ;
 wire \top_I.branch[1].l_um_ena[14] ;
 wire \top_I.branch[1].l_um_ena[15] ;
 wire \top_I.branch[1].l_um_ena[1] ;
 wire \top_I.branch[1].l_um_ena[2] ;
 wire \top_I.branch[1].l_um_ena[3] ;
 wire \top_I.branch[1].l_um_ena[4] ;
 wire \top_I.branch[1].l_um_ena[5] ;
 wire \top_I.branch[1].l_um_ena[6] ;
 wire \top_I.branch[1].l_um_ena[7] ;
 wire \top_I.branch[1].l_um_ena[8] ;
 wire \top_I.branch[1].l_um_ena[9] ;
 wire \top_I.branch[1].l_um_iw[0] ;
 wire \top_I.branch[1].l_um_iw[100] ;
 wire \top_I.branch[1].l_um_iw[101] ;
 wire \top_I.branch[1].l_um_iw[102] ;
 wire \top_I.branch[1].l_um_iw[103] ;
 wire \top_I.branch[1].l_um_iw[104] ;
 wire \top_I.branch[1].l_um_iw[105] ;
 wire \top_I.branch[1].l_um_iw[106] ;
 wire \top_I.branch[1].l_um_iw[107] ;
 wire \top_I.branch[1].l_um_iw[108] ;
 wire \top_I.branch[1].l_um_iw[109] ;
 wire \top_I.branch[1].l_um_iw[10] ;
 wire \top_I.branch[1].l_um_iw[110] ;
 wire \top_I.branch[1].l_um_iw[111] ;
 wire \top_I.branch[1].l_um_iw[112] ;
 wire \top_I.branch[1].l_um_iw[113] ;
 wire \top_I.branch[1].l_um_iw[114] ;
 wire \top_I.branch[1].l_um_iw[115] ;
 wire \top_I.branch[1].l_um_iw[116] ;
 wire \top_I.branch[1].l_um_iw[117] ;
 wire \top_I.branch[1].l_um_iw[118] ;
 wire \top_I.branch[1].l_um_iw[119] ;
 wire \top_I.branch[1].l_um_iw[11] ;
 wire \top_I.branch[1].l_um_iw[120] ;
 wire \top_I.branch[1].l_um_iw[121] ;
 wire \top_I.branch[1].l_um_iw[122] ;
 wire \top_I.branch[1].l_um_iw[123] ;
 wire \top_I.branch[1].l_um_iw[124] ;
 wire \top_I.branch[1].l_um_iw[125] ;
 wire \top_I.branch[1].l_um_iw[126] ;
 wire \top_I.branch[1].l_um_iw[127] ;
 wire \top_I.branch[1].l_um_iw[128] ;
 wire \top_I.branch[1].l_um_iw[129] ;
 wire \top_I.branch[1].l_um_iw[12] ;
 wire \top_I.branch[1].l_um_iw[130] ;
 wire \top_I.branch[1].l_um_iw[131] ;
 wire \top_I.branch[1].l_um_iw[132] ;
 wire \top_I.branch[1].l_um_iw[133] ;
 wire \top_I.branch[1].l_um_iw[134] ;
 wire \top_I.branch[1].l_um_iw[135] ;
 wire \top_I.branch[1].l_um_iw[136] ;
 wire \top_I.branch[1].l_um_iw[137] ;
 wire \top_I.branch[1].l_um_iw[138] ;
 wire \top_I.branch[1].l_um_iw[139] ;
 wire \top_I.branch[1].l_um_iw[13] ;
 wire \top_I.branch[1].l_um_iw[140] ;
 wire \top_I.branch[1].l_um_iw[141] ;
 wire \top_I.branch[1].l_um_iw[142] ;
 wire \top_I.branch[1].l_um_iw[143] ;
 wire \top_I.branch[1].l_um_iw[144] ;
 wire \top_I.branch[1].l_um_iw[145] ;
 wire \top_I.branch[1].l_um_iw[146] ;
 wire \top_I.branch[1].l_um_iw[147] ;
 wire \top_I.branch[1].l_um_iw[148] ;
 wire \top_I.branch[1].l_um_iw[149] ;
 wire \top_I.branch[1].l_um_iw[14] ;
 wire \top_I.branch[1].l_um_iw[150] ;
 wire \top_I.branch[1].l_um_iw[151] ;
 wire \top_I.branch[1].l_um_iw[152] ;
 wire \top_I.branch[1].l_um_iw[153] ;
 wire \top_I.branch[1].l_um_iw[154] ;
 wire \top_I.branch[1].l_um_iw[155] ;
 wire \top_I.branch[1].l_um_iw[156] ;
 wire \top_I.branch[1].l_um_iw[157] ;
 wire \top_I.branch[1].l_um_iw[158] ;
 wire \top_I.branch[1].l_um_iw[159] ;
 wire \top_I.branch[1].l_um_iw[15] ;
 wire \top_I.branch[1].l_um_iw[160] ;
 wire \top_I.branch[1].l_um_iw[161] ;
 wire \top_I.branch[1].l_um_iw[162] ;
 wire \top_I.branch[1].l_um_iw[163] ;
 wire \top_I.branch[1].l_um_iw[164] ;
 wire \top_I.branch[1].l_um_iw[165] ;
 wire \top_I.branch[1].l_um_iw[166] ;
 wire \top_I.branch[1].l_um_iw[167] ;
 wire \top_I.branch[1].l_um_iw[168] ;
 wire \top_I.branch[1].l_um_iw[169] ;
 wire \top_I.branch[1].l_um_iw[16] ;
 wire \top_I.branch[1].l_um_iw[170] ;
 wire \top_I.branch[1].l_um_iw[171] ;
 wire \top_I.branch[1].l_um_iw[172] ;
 wire \top_I.branch[1].l_um_iw[173] ;
 wire \top_I.branch[1].l_um_iw[174] ;
 wire \top_I.branch[1].l_um_iw[175] ;
 wire \top_I.branch[1].l_um_iw[176] ;
 wire \top_I.branch[1].l_um_iw[177] ;
 wire \top_I.branch[1].l_um_iw[178] ;
 wire \top_I.branch[1].l_um_iw[179] ;
 wire \top_I.branch[1].l_um_iw[17] ;
 wire \top_I.branch[1].l_um_iw[180] ;
 wire \top_I.branch[1].l_um_iw[181] ;
 wire \top_I.branch[1].l_um_iw[182] ;
 wire \top_I.branch[1].l_um_iw[183] ;
 wire \top_I.branch[1].l_um_iw[184] ;
 wire \top_I.branch[1].l_um_iw[185] ;
 wire \top_I.branch[1].l_um_iw[186] ;
 wire \top_I.branch[1].l_um_iw[187] ;
 wire \top_I.branch[1].l_um_iw[188] ;
 wire \top_I.branch[1].l_um_iw[189] ;
 wire \top_I.branch[1].l_um_iw[18] ;
 wire \top_I.branch[1].l_um_iw[190] ;
 wire \top_I.branch[1].l_um_iw[191] ;
 wire \top_I.branch[1].l_um_iw[192] ;
 wire \top_I.branch[1].l_um_iw[193] ;
 wire \top_I.branch[1].l_um_iw[194] ;
 wire \top_I.branch[1].l_um_iw[195] ;
 wire \top_I.branch[1].l_um_iw[196] ;
 wire \top_I.branch[1].l_um_iw[197] ;
 wire \top_I.branch[1].l_um_iw[198] ;
 wire \top_I.branch[1].l_um_iw[199] ;
 wire \top_I.branch[1].l_um_iw[19] ;
 wire \top_I.branch[1].l_um_iw[1] ;
 wire \top_I.branch[1].l_um_iw[200] ;
 wire \top_I.branch[1].l_um_iw[201] ;
 wire \top_I.branch[1].l_um_iw[202] ;
 wire \top_I.branch[1].l_um_iw[203] ;
 wire \top_I.branch[1].l_um_iw[204] ;
 wire \top_I.branch[1].l_um_iw[205] ;
 wire \top_I.branch[1].l_um_iw[206] ;
 wire \top_I.branch[1].l_um_iw[207] ;
 wire \top_I.branch[1].l_um_iw[208] ;
 wire \top_I.branch[1].l_um_iw[209] ;
 wire \top_I.branch[1].l_um_iw[20] ;
 wire \top_I.branch[1].l_um_iw[210] ;
 wire \top_I.branch[1].l_um_iw[211] ;
 wire \top_I.branch[1].l_um_iw[212] ;
 wire \top_I.branch[1].l_um_iw[213] ;
 wire \top_I.branch[1].l_um_iw[214] ;
 wire \top_I.branch[1].l_um_iw[215] ;
 wire \top_I.branch[1].l_um_iw[216] ;
 wire \top_I.branch[1].l_um_iw[217] ;
 wire \top_I.branch[1].l_um_iw[218] ;
 wire \top_I.branch[1].l_um_iw[219] ;
 wire \top_I.branch[1].l_um_iw[21] ;
 wire \top_I.branch[1].l_um_iw[220] ;
 wire \top_I.branch[1].l_um_iw[221] ;
 wire \top_I.branch[1].l_um_iw[222] ;
 wire \top_I.branch[1].l_um_iw[223] ;
 wire \top_I.branch[1].l_um_iw[224] ;
 wire \top_I.branch[1].l_um_iw[225] ;
 wire \top_I.branch[1].l_um_iw[226] ;
 wire \top_I.branch[1].l_um_iw[227] ;
 wire \top_I.branch[1].l_um_iw[228] ;
 wire \top_I.branch[1].l_um_iw[229] ;
 wire \top_I.branch[1].l_um_iw[22] ;
 wire \top_I.branch[1].l_um_iw[230] ;
 wire \top_I.branch[1].l_um_iw[231] ;
 wire \top_I.branch[1].l_um_iw[232] ;
 wire \top_I.branch[1].l_um_iw[233] ;
 wire \top_I.branch[1].l_um_iw[234] ;
 wire \top_I.branch[1].l_um_iw[235] ;
 wire \top_I.branch[1].l_um_iw[236] ;
 wire \top_I.branch[1].l_um_iw[237] ;
 wire \top_I.branch[1].l_um_iw[238] ;
 wire \top_I.branch[1].l_um_iw[239] ;
 wire \top_I.branch[1].l_um_iw[23] ;
 wire \top_I.branch[1].l_um_iw[240] ;
 wire \top_I.branch[1].l_um_iw[241] ;
 wire \top_I.branch[1].l_um_iw[242] ;
 wire \top_I.branch[1].l_um_iw[243] ;
 wire \top_I.branch[1].l_um_iw[244] ;
 wire \top_I.branch[1].l_um_iw[245] ;
 wire \top_I.branch[1].l_um_iw[246] ;
 wire \top_I.branch[1].l_um_iw[247] ;
 wire \top_I.branch[1].l_um_iw[248] ;
 wire \top_I.branch[1].l_um_iw[249] ;
 wire \top_I.branch[1].l_um_iw[24] ;
 wire \top_I.branch[1].l_um_iw[250] ;
 wire \top_I.branch[1].l_um_iw[251] ;
 wire \top_I.branch[1].l_um_iw[252] ;
 wire \top_I.branch[1].l_um_iw[253] ;
 wire \top_I.branch[1].l_um_iw[254] ;
 wire \top_I.branch[1].l_um_iw[255] ;
 wire \top_I.branch[1].l_um_iw[256] ;
 wire \top_I.branch[1].l_um_iw[257] ;
 wire \top_I.branch[1].l_um_iw[258] ;
 wire \top_I.branch[1].l_um_iw[259] ;
 wire \top_I.branch[1].l_um_iw[25] ;
 wire \top_I.branch[1].l_um_iw[260] ;
 wire \top_I.branch[1].l_um_iw[261] ;
 wire \top_I.branch[1].l_um_iw[262] ;
 wire \top_I.branch[1].l_um_iw[263] ;
 wire \top_I.branch[1].l_um_iw[264] ;
 wire \top_I.branch[1].l_um_iw[265] ;
 wire \top_I.branch[1].l_um_iw[266] ;
 wire \top_I.branch[1].l_um_iw[267] ;
 wire \top_I.branch[1].l_um_iw[268] ;
 wire \top_I.branch[1].l_um_iw[269] ;
 wire \top_I.branch[1].l_um_iw[26] ;
 wire \top_I.branch[1].l_um_iw[270] ;
 wire \top_I.branch[1].l_um_iw[271] ;
 wire \top_I.branch[1].l_um_iw[272] ;
 wire \top_I.branch[1].l_um_iw[273] ;
 wire \top_I.branch[1].l_um_iw[274] ;
 wire \top_I.branch[1].l_um_iw[275] ;
 wire \top_I.branch[1].l_um_iw[276] ;
 wire \top_I.branch[1].l_um_iw[277] ;
 wire \top_I.branch[1].l_um_iw[278] ;
 wire \top_I.branch[1].l_um_iw[279] ;
 wire \top_I.branch[1].l_um_iw[27] ;
 wire \top_I.branch[1].l_um_iw[280] ;
 wire \top_I.branch[1].l_um_iw[281] ;
 wire \top_I.branch[1].l_um_iw[282] ;
 wire \top_I.branch[1].l_um_iw[283] ;
 wire \top_I.branch[1].l_um_iw[284] ;
 wire \top_I.branch[1].l_um_iw[285] ;
 wire \top_I.branch[1].l_um_iw[286] ;
 wire \top_I.branch[1].l_um_iw[287] ;
 wire \top_I.branch[1].l_um_iw[28] ;
 wire \top_I.branch[1].l_um_iw[29] ;
 wire \top_I.branch[1].l_um_iw[2] ;
 wire \top_I.branch[1].l_um_iw[30] ;
 wire \top_I.branch[1].l_um_iw[31] ;
 wire \top_I.branch[1].l_um_iw[32] ;
 wire \top_I.branch[1].l_um_iw[33] ;
 wire \top_I.branch[1].l_um_iw[34] ;
 wire \top_I.branch[1].l_um_iw[35] ;
 wire \top_I.branch[1].l_um_iw[36] ;
 wire \top_I.branch[1].l_um_iw[37] ;
 wire \top_I.branch[1].l_um_iw[38] ;
 wire \top_I.branch[1].l_um_iw[39] ;
 wire \top_I.branch[1].l_um_iw[3] ;
 wire \top_I.branch[1].l_um_iw[40] ;
 wire \top_I.branch[1].l_um_iw[41] ;
 wire \top_I.branch[1].l_um_iw[42] ;
 wire \top_I.branch[1].l_um_iw[43] ;
 wire \top_I.branch[1].l_um_iw[44] ;
 wire \top_I.branch[1].l_um_iw[45] ;
 wire \top_I.branch[1].l_um_iw[46] ;
 wire \top_I.branch[1].l_um_iw[47] ;
 wire \top_I.branch[1].l_um_iw[48] ;
 wire \top_I.branch[1].l_um_iw[49] ;
 wire \top_I.branch[1].l_um_iw[4] ;
 wire \top_I.branch[1].l_um_iw[50] ;
 wire \top_I.branch[1].l_um_iw[51] ;
 wire \top_I.branch[1].l_um_iw[52] ;
 wire \top_I.branch[1].l_um_iw[53] ;
 wire \top_I.branch[1].l_um_iw[54] ;
 wire \top_I.branch[1].l_um_iw[55] ;
 wire \top_I.branch[1].l_um_iw[56] ;
 wire \top_I.branch[1].l_um_iw[57] ;
 wire \top_I.branch[1].l_um_iw[58] ;
 wire \top_I.branch[1].l_um_iw[59] ;
 wire \top_I.branch[1].l_um_iw[5] ;
 wire \top_I.branch[1].l_um_iw[60] ;
 wire \top_I.branch[1].l_um_iw[61] ;
 wire \top_I.branch[1].l_um_iw[62] ;
 wire \top_I.branch[1].l_um_iw[63] ;
 wire \top_I.branch[1].l_um_iw[64] ;
 wire \top_I.branch[1].l_um_iw[65] ;
 wire \top_I.branch[1].l_um_iw[66] ;
 wire \top_I.branch[1].l_um_iw[67] ;
 wire \top_I.branch[1].l_um_iw[68] ;
 wire \top_I.branch[1].l_um_iw[69] ;
 wire \top_I.branch[1].l_um_iw[6] ;
 wire \top_I.branch[1].l_um_iw[70] ;
 wire \top_I.branch[1].l_um_iw[71] ;
 wire \top_I.branch[1].l_um_iw[72] ;
 wire \top_I.branch[1].l_um_iw[73] ;
 wire \top_I.branch[1].l_um_iw[74] ;
 wire \top_I.branch[1].l_um_iw[75] ;
 wire \top_I.branch[1].l_um_iw[76] ;
 wire \top_I.branch[1].l_um_iw[77] ;
 wire \top_I.branch[1].l_um_iw[78] ;
 wire \top_I.branch[1].l_um_iw[79] ;
 wire \top_I.branch[1].l_um_iw[7] ;
 wire \top_I.branch[1].l_um_iw[80] ;
 wire \top_I.branch[1].l_um_iw[81] ;
 wire \top_I.branch[1].l_um_iw[82] ;
 wire \top_I.branch[1].l_um_iw[83] ;
 wire \top_I.branch[1].l_um_iw[84] ;
 wire \top_I.branch[1].l_um_iw[85] ;
 wire \top_I.branch[1].l_um_iw[86] ;
 wire \top_I.branch[1].l_um_iw[87] ;
 wire \top_I.branch[1].l_um_iw[88] ;
 wire \top_I.branch[1].l_um_iw[89] ;
 wire \top_I.branch[1].l_um_iw[8] ;
 wire \top_I.branch[1].l_um_iw[90] ;
 wire \top_I.branch[1].l_um_iw[91] ;
 wire \top_I.branch[1].l_um_iw[92] ;
 wire \top_I.branch[1].l_um_iw[93] ;
 wire \top_I.branch[1].l_um_iw[94] ;
 wire \top_I.branch[1].l_um_iw[95] ;
 wire \top_I.branch[1].l_um_iw[96] ;
 wire \top_I.branch[1].l_um_iw[97] ;
 wire \top_I.branch[1].l_um_iw[98] ;
 wire \top_I.branch[1].l_um_iw[99] ;
 wire \top_I.branch[1].l_um_iw[9] ;
 wire \top_I.branch[1].l_um_k_zero[0] ;
 wire \top_I.branch[1].l_um_k_zero[10] ;
 wire \top_I.branch[1].l_um_k_zero[11] ;
 wire \top_I.branch[1].l_um_k_zero[12] ;
 wire \top_I.branch[1].l_um_k_zero[13] ;
 wire \top_I.branch[1].l_um_k_zero[14] ;
 wire \top_I.branch[1].l_um_k_zero[15] ;
 wire \top_I.branch[1].l_um_k_zero[1] ;
 wire \top_I.branch[1].l_um_k_zero[2] ;
 wire \top_I.branch[1].l_um_k_zero[3] ;
 wire \top_I.branch[1].l_um_k_zero[4] ;
 wire \top_I.branch[1].l_um_k_zero[5] ;
 wire \top_I.branch[1].l_um_k_zero[6] ;
 wire \top_I.branch[1].l_um_k_zero[7] ;
 wire \top_I.branch[1].l_um_k_zero[8] ;
 wire \top_I.branch[1].l_um_k_zero[9] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[20].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[20].l_k_one ;
 wire \top_I.branch[20].l_k_zero ;
 wire \top_I.branch[20].l_um_ena[0] ;
 wire \top_I.branch[20].l_um_ena[10] ;
 wire \top_I.branch[20].l_um_ena[11] ;
 wire \top_I.branch[20].l_um_ena[12] ;
 wire \top_I.branch[20].l_um_ena[13] ;
 wire \top_I.branch[20].l_um_ena[14] ;
 wire \top_I.branch[20].l_um_ena[15] ;
 wire \top_I.branch[20].l_um_ena[1] ;
 wire \top_I.branch[20].l_um_ena[2] ;
 wire \top_I.branch[20].l_um_ena[3] ;
 wire \top_I.branch[20].l_um_ena[4] ;
 wire \top_I.branch[20].l_um_ena[5] ;
 wire \top_I.branch[20].l_um_ena[6] ;
 wire \top_I.branch[20].l_um_ena[7] ;
 wire \top_I.branch[20].l_um_ena[8] ;
 wire \top_I.branch[20].l_um_ena[9] ;
 wire \top_I.branch[20].l_um_iw[0] ;
 wire \top_I.branch[20].l_um_iw[100] ;
 wire \top_I.branch[20].l_um_iw[101] ;
 wire \top_I.branch[20].l_um_iw[102] ;
 wire \top_I.branch[20].l_um_iw[103] ;
 wire \top_I.branch[20].l_um_iw[104] ;
 wire \top_I.branch[20].l_um_iw[105] ;
 wire \top_I.branch[20].l_um_iw[106] ;
 wire \top_I.branch[20].l_um_iw[107] ;
 wire \top_I.branch[20].l_um_iw[108] ;
 wire \top_I.branch[20].l_um_iw[109] ;
 wire \top_I.branch[20].l_um_iw[10] ;
 wire \top_I.branch[20].l_um_iw[110] ;
 wire \top_I.branch[20].l_um_iw[111] ;
 wire \top_I.branch[20].l_um_iw[112] ;
 wire \top_I.branch[20].l_um_iw[113] ;
 wire \top_I.branch[20].l_um_iw[114] ;
 wire \top_I.branch[20].l_um_iw[115] ;
 wire \top_I.branch[20].l_um_iw[116] ;
 wire \top_I.branch[20].l_um_iw[117] ;
 wire \top_I.branch[20].l_um_iw[118] ;
 wire \top_I.branch[20].l_um_iw[119] ;
 wire \top_I.branch[20].l_um_iw[11] ;
 wire \top_I.branch[20].l_um_iw[120] ;
 wire \top_I.branch[20].l_um_iw[121] ;
 wire \top_I.branch[20].l_um_iw[122] ;
 wire \top_I.branch[20].l_um_iw[123] ;
 wire \top_I.branch[20].l_um_iw[124] ;
 wire \top_I.branch[20].l_um_iw[125] ;
 wire \top_I.branch[20].l_um_iw[126] ;
 wire \top_I.branch[20].l_um_iw[127] ;
 wire \top_I.branch[20].l_um_iw[128] ;
 wire \top_I.branch[20].l_um_iw[129] ;
 wire \top_I.branch[20].l_um_iw[12] ;
 wire \top_I.branch[20].l_um_iw[130] ;
 wire \top_I.branch[20].l_um_iw[131] ;
 wire \top_I.branch[20].l_um_iw[132] ;
 wire \top_I.branch[20].l_um_iw[133] ;
 wire \top_I.branch[20].l_um_iw[134] ;
 wire \top_I.branch[20].l_um_iw[135] ;
 wire \top_I.branch[20].l_um_iw[136] ;
 wire \top_I.branch[20].l_um_iw[137] ;
 wire \top_I.branch[20].l_um_iw[138] ;
 wire \top_I.branch[20].l_um_iw[139] ;
 wire \top_I.branch[20].l_um_iw[13] ;
 wire \top_I.branch[20].l_um_iw[140] ;
 wire \top_I.branch[20].l_um_iw[141] ;
 wire \top_I.branch[20].l_um_iw[142] ;
 wire \top_I.branch[20].l_um_iw[143] ;
 wire \top_I.branch[20].l_um_iw[144] ;
 wire \top_I.branch[20].l_um_iw[145] ;
 wire \top_I.branch[20].l_um_iw[146] ;
 wire \top_I.branch[20].l_um_iw[147] ;
 wire \top_I.branch[20].l_um_iw[148] ;
 wire \top_I.branch[20].l_um_iw[149] ;
 wire \top_I.branch[20].l_um_iw[14] ;
 wire \top_I.branch[20].l_um_iw[150] ;
 wire \top_I.branch[20].l_um_iw[151] ;
 wire \top_I.branch[20].l_um_iw[152] ;
 wire \top_I.branch[20].l_um_iw[153] ;
 wire \top_I.branch[20].l_um_iw[154] ;
 wire \top_I.branch[20].l_um_iw[155] ;
 wire \top_I.branch[20].l_um_iw[156] ;
 wire \top_I.branch[20].l_um_iw[157] ;
 wire \top_I.branch[20].l_um_iw[158] ;
 wire \top_I.branch[20].l_um_iw[159] ;
 wire \top_I.branch[20].l_um_iw[15] ;
 wire \top_I.branch[20].l_um_iw[160] ;
 wire \top_I.branch[20].l_um_iw[161] ;
 wire \top_I.branch[20].l_um_iw[162] ;
 wire \top_I.branch[20].l_um_iw[163] ;
 wire \top_I.branch[20].l_um_iw[164] ;
 wire \top_I.branch[20].l_um_iw[165] ;
 wire \top_I.branch[20].l_um_iw[166] ;
 wire \top_I.branch[20].l_um_iw[167] ;
 wire \top_I.branch[20].l_um_iw[168] ;
 wire \top_I.branch[20].l_um_iw[169] ;
 wire \top_I.branch[20].l_um_iw[16] ;
 wire \top_I.branch[20].l_um_iw[170] ;
 wire \top_I.branch[20].l_um_iw[171] ;
 wire \top_I.branch[20].l_um_iw[172] ;
 wire \top_I.branch[20].l_um_iw[173] ;
 wire \top_I.branch[20].l_um_iw[174] ;
 wire \top_I.branch[20].l_um_iw[175] ;
 wire \top_I.branch[20].l_um_iw[176] ;
 wire \top_I.branch[20].l_um_iw[177] ;
 wire \top_I.branch[20].l_um_iw[178] ;
 wire \top_I.branch[20].l_um_iw[179] ;
 wire \top_I.branch[20].l_um_iw[17] ;
 wire \top_I.branch[20].l_um_iw[180] ;
 wire \top_I.branch[20].l_um_iw[181] ;
 wire \top_I.branch[20].l_um_iw[182] ;
 wire \top_I.branch[20].l_um_iw[183] ;
 wire \top_I.branch[20].l_um_iw[184] ;
 wire \top_I.branch[20].l_um_iw[185] ;
 wire \top_I.branch[20].l_um_iw[186] ;
 wire \top_I.branch[20].l_um_iw[187] ;
 wire \top_I.branch[20].l_um_iw[188] ;
 wire \top_I.branch[20].l_um_iw[189] ;
 wire \top_I.branch[20].l_um_iw[18] ;
 wire \top_I.branch[20].l_um_iw[190] ;
 wire \top_I.branch[20].l_um_iw[191] ;
 wire \top_I.branch[20].l_um_iw[192] ;
 wire \top_I.branch[20].l_um_iw[193] ;
 wire \top_I.branch[20].l_um_iw[194] ;
 wire \top_I.branch[20].l_um_iw[195] ;
 wire \top_I.branch[20].l_um_iw[196] ;
 wire \top_I.branch[20].l_um_iw[197] ;
 wire \top_I.branch[20].l_um_iw[198] ;
 wire \top_I.branch[20].l_um_iw[199] ;
 wire \top_I.branch[20].l_um_iw[19] ;
 wire \top_I.branch[20].l_um_iw[1] ;
 wire \top_I.branch[20].l_um_iw[200] ;
 wire \top_I.branch[20].l_um_iw[201] ;
 wire \top_I.branch[20].l_um_iw[202] ;
 wire \top_I.branch[20].l_um_iw[203] ;
 wire \top_I.branch[20].l_um_iw[204] ;
 wire \top_I.branch[20].l_um_iw[205] ;
 wire \top_I.branch[20].l_um_iw[206] ;
 wire \top_I.branch[20].l_um_iw[207] ;
 wire \top_I.branch[20].l_um_iw[208] ;
 wire \top_I.branch[20].l_um_iw[209] ;
 wire \top_I.branch[20].l_um_iw[20] ;
 wire \top_I.branch[20].l_um_iw[210] ;
 wire \top_I.branch[20].l_um_iw[211] ;
 wire \top_I.branch[20].l_um_iw[212] ;
 wire \top_I.branch[20].l_um_iw[213] ;
 wire \top_I.branch[20].l_um_iw[214] ;
 wire \top_I.branch[20].l_um_iw[215] ;
 wire \top_I.branch[20].l_um_iw[216] ;
 wire \top_I.branch[20].l_um_iw[217] ;
 wire \top_I.branch[20].l_um_iw[218] ;
 wire \top_I.branch[20].l_um_iw[219] ;
 wire \top_I.branch[20].l_um_iw[21] ;
 wire \top_I.branch[20].l_um_iw[220] ;
 wire \top_I.branch[20].l_um_iw[221] ;
 wire \top_I.branch[20].l_um_iw[222] ;
 wire \top_I.branch[20].l_um_iw[223] ;
 wire \top_I.branch[20].l_um_iw[224] ;
 wire \top_I.branch[20].l_um_iw[225] ;
 wire \top_I.branch[20].l_um_iw[226] ;
 wire \top_I.branch[20].l_um_iw[227] ;
 wire \top_I.branch[20].l_um_iw[228] ;
 wire \top_I.branch[20].l_um_iw[229] ;
 wire \top_I.branch[20].l_um_iw[22] ;
 wire \top_I.branch[20].l_um_iw[230] ;
 wire \top_I.branch[20].l_um_iw[231] ;
 wire \top_I.branch[20].l_um_iw[232] ;
 wire \top_I.branch[20].l_um_iw[233] ;
 wire \top_I.branch[20].l_um_iw[234] ;
 wire \top_I.branch[20].l_um_iw[235] ;
 wire \top_I.branch[20].l_um_iw[236] ;
 wire \top_I.branch[20].l_um_iw[237] ;
 wire \top_I.branch[20].l_um_iw[238] ;
 wire \top_I.branch[20].l_um_iw[239] ;
 wire \top_I.branch[20].l_um_iw[23] ;
 wire \top_I.branch[20].l_um_iw[240] ;
 wire \top_I.branch[20].l_um_iw[241] ;
 wire \top_I.branch[20].l_um_iw[242] ;
 wire \top_I.branch[20].l_um_iw[243] ;
 wire \top_I.branch[20].l_um_iw[244] ;
 wire \top_I.branch[20].l_um_iw[245] ;
 wire \top_I.branch[20].l_um_iw[246] ;
 wire \top_I.branch[20].l_um_iw[247] ;
 wire \top_I.branch[20].l_um_iw[248] ;
 wire \top_I.branch[20].l_um_iw[249] ;
 wire \top_I.branch[20].l_um_iw[24] ;
 wire \top_I.branch[20].l_um_iw[250] ;
 wire \top_I.branch[20].l_um_iw[251] ;
 wire \top_I.branch[20].l_um_iw[252] ;
 wire \top_I.branch[20].l_um_iw[253] ;
 wire \top_I.branch[20].l_um_iw[254] ;
 wire \top_I.branch[20].l_um_iw[255] ;
 wire \top_I.branch[20].l_um_iw[256] ;
 wire \top_I.branch[20].l_um_iw[257] ;
 wire \top_I.branch[20].l_um_iw[258] ;
 wire \top_I.branch[20].l_um_iw[259] ;
 wire \top_I.branch[20].l_um_iw[25] ;
 wire \top_I.branch[20].l_um_iw[260] ;
 wire \top_I.branch[20].l_um_iw[261] ;
 wire \top_I.branch[20].l_um_iw[262] ;
 wire \top_I.branch[20].l_um_iw[263] ;
 wire \top_I.branch[20].l_um_iw[264] ;
 wire \top_I.branch[20].l_um_iw[265] ;
 wire \top_I.branch[20].l_um_iw[266] ;
 wire \top_I.branch[20].l_um_iw[267] ;
 wire \top_I.branch[20].l_um_iw[268] ;
 wire \top_I.branch[20].l_um_iw[269] ;
 wire \top_I.branch[20].l_um_iw[26] ;
 wire \top_I.branch[20].l_um_iw[270] ;
 wire \top_I.branch[20].l_um_iw[271] ;
 wire \top_I.branch[20].l_um_iw[272] ;
 wire \top_I.branch[20].l_um_iw[273] ;
 wire \top_I.branch[20].l_um_iw[274] ;
 wire \top_I.branch[20].l_um_iw[275] ;
 wire \top_I.branch[20].l_um_iw[276] ;
 wire \top_I.branch[20].l_um_iw[277] ;
 wire \top_I.branch[20].l_um_iw[278] ;
 wire \top_I.branch[20].l_um_iw[279] ;
 wire \top_I.branch[20].l_um_iw[27] ;
 wire \top_I.branch[20].l_um_iw[280] ;
 wire \top_I.branch[20].l_um_iw[281] ;
 wire \top_I.branch[20].l_um_iw[282] ;
 wire \top_I.branch[20].l_um_iw[283] ;
 wire \top_I.branch[20].l_um_iw[284] ;
 wire \top_I.branch[20].l_um_iw[285] ;
 wire \top_I.branch[20].l_um_iw[286] ;
 wire \top_I.branch[20].l_um_iw[287] ;
 wire \top_I.branch[20].l_um_iw[28] ;
 wire \top_I.branch[20].l_um_iw[29] ;
 wire \top_I.branch[20].l_um_iw[2] ;
 wire \top_I.branch[20].l_um_iw[30] ;
 wire \top_I.branch[20].l_um_iw[31] ;
 wire \top_I.branch[20].l_um_iw[32] ;
 wire \top_I.branch[20].l_um_iw[33] ;
 wire \top_I.branch[20].l_um_iw[34] ;
 wire \top_I.branch[20].l_um_iw[35] ;
 wire \top_I.branch[20].l_um_iw[36] ;
 wire \top_I.branch[20].l_um_iw[37] ;
 wire \top_I.branch[20].l_um_iw[38] ;
 wire \top_I.branch[20].l_um_iw[39] ;
 wire \top_I.branch[20].l_um_iw[3] ;
 wire \top_I.branch[20].l_um_iw[40] ;
 wire \top_I.branch[20].l_um_iw[41] ;
 wire \top_I.branch[20].l_um_iw[42] ;
 wire \top_I.branch[20].l_um_iw[43] ;
 wire \top_I.branch[20].l_um_iw[44] ;
 wire \top_I.branch[20].l_um_iw[45] ;
 wire \top_I.branch[20].l_um_iw[46] ;
 wire \top_I.branch[20].l_um_iw[47] ;
 wire \top_I.branch[20].l_um_iw[48] ;
 wire \top_I.branch[20].l_um_iw[49] ;
 wire \top_I.branch[20].l_um_iw[4] ;
 wire \top_I.branch[20].l_um_iw[50] ;
 wire \top_I.branch[20].l_um_iw[51] ;
 wire \top_I.branch[20].l_um_iw[52] ;
 wire \top_I.branch[20].l_um_iw[53] ;
 wire \top_I.branch[20].l_um_iw[54] ;
 wire \top_I.branch[20].l_um_iw[55] ;
 wire \top_I.branch[20].l_um_iw[56] ;
 wire \top_I.branch[20].l_um_iw[57] ;
 wire \top_I.branch[20].l_um_iw[58] ;
 wire \top_I.branch[20].l_um_iw[59] ;
 wire \top_I.branch[20].l_um_iw[5] ;
 wire \top_I.branch[20].l_um_iw[60] ;
 wire \top_I.branch[20].l_um_iw[61] ;
 wire \top_I.branch[20].l_um_iw[62] ;
 wire \top_I.branch[20].l_um_iw[63] ;
 wire \top_I.branch[20].l_um_iw[64] ;
 wire \top_I.branch[20].l_um_iw[65] ;
 wire \top_I.branch[20].l_um_iw[66] ;
 wire \top_I.branch[20].l_um_iw[67] ;
 wire \top_I.branch[20].l_um_iw[68] ;
 wire \top_I.branch[20].l_um_iw[69] ;
 wire \top_I.branch[20].l_um_iw[6] ;
 wire \top_I.branch[20].l_um_iw[70] ;
 wire \top_I.branch[20].l_um_iw[71] ;
 wire \top_I.branch[20].l_um_iw[72] ;
 wire \top_I.branch[20].l_um_iw[73] ;
 wire \top_I.branch[20].l_um_iw[74] ;
 wire \top_I.branch[20].l_um_iw[75] ;
 wire \top_I.branch[20].l_um_iw[76] ;
 wire \top_I.branch[20].l_um_iw[77] ;
 wire \top_I.branch[20].l_um_iw[78] ;
 wire \top_I.branch[20].l_um_iw[79] ;
 wire \top_I.branch[20].l_um_iw[7] ;
 wire \top_I.branch[20].l_um_iw[80] ;
 wire \top_I.branch[20].l_um_iw[81] ;
 wire \top_I.branch[20].l_um_iw[82] ;
 wire \top_I.branch[20].l_um_iw[83] ;
 wire \top_I.branch[20].l_um_iw[84] ;
 wire \top_I.branch[20].l_um_iw[85] ;
 wire \top_I.branch[20].l_um_iw[86] ;
 wire \top_I.branch[20].l_um_iw[87] ;
 wire \top_I.branch[20].l_um_iw[88] ;
 wire \top_I.branch[20].l_um_iw[89] ;
 wire \top_I.branch[20].l_um_iw[8] ;
 wire \top_I.branch[20].l_um_iw[90] ;
 wire \top_I.branch[20].l_um_iw[91] ;
 wire \top_I.branch[20].l_um_iw[92] ;
 wire \top_I.branch[20].l_um_iw[93] ;
 wire \top_I.branch[20].l_um_iw[94] ;
 wire \top_I.branch[20].l_um_iw[95] ;
 wire \top_I.branch[20].l_um_iw[96] ;
 wire \top_I.branch[20].l_um_iw[97] ;
 wire \top_I.branch[20].l_um_iw[98] ;
 wire \top_I.branch[20].l_um_iw[99] ;
 wire \top_I.branch[20].l_um_iw[9] ;
 wire \top_I.branch[20].l_um_k_zero[0] ;
 wire \top_I.branch[20].l_um_k_zero[10] ;
 wire \top_I.branch[20].l_um_k_zero[11] ;
 wire \top_I.branch[20].l_um_k_zero[12] ;
 wire \top_I.branch[20].l_um_k_zero[13] ;
 wire \top_I.branch[20].l_um_k_zero[14] ;
 wire \top_I.branch[20].l_um_k_zero[15] ;
 wire \top_I.branch[20].l_um_k_zero[1] ;
 wire \top_I.branch[20].l_um_k_zero[2] ;
 wire \top_I.branch[20].l_um_k_zero[3] ;
 wire \top_I.branch[20].l_um_k_zero[4] ;
 wire \top_I.branch[20].l_um_k_zero[5] ;
 wire \top_I.branch[20].l_um_k_zero[6] ;
 wire \top_I.branch[20].l_um_k_zero[7] ;
 wire \top_I.branch[20].l_um_k_zero[8] ;
 wire \top_I.branch[20].l_um_k_zero[9] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[21].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[21].l_k_one ;
 wire \top_I.branch[21].l_k_zero ;
 wire \top_I.branch[21].l_um_ena[0] ;
 wire \top_I.branch[21].l_um_ena[10] ;
 wire \top_I.branch[21].l_um_ena[11] ;
 wire \top_I.branch[21].l_um_ena[12] ;
 wire \top_I.branch[21].l_um_ena[13] ;
 wire \top_I.branch[21].l_um_ena[14] ;
 wire \top_I.branch[21].l_um_ena[15] ;
 wire \top_I.branch[21].l_um_ena[1] ;
 wire \top_I.branch[21].l_um_ena[2] ;
 wire \top_I.branch[21].l_um_ena[3] ;
 wire \top_I.branch[21].l_um_ena[4] ;
 wire \top_I.branch[21].l_um_ena[5] ;
 wire \top_I.branch[21].l_um_ena[6] ;
 wire \top_I.branch[21].l_um_ena[7] ;
 wire \top_I.branch[21].l_um_ena[8] ;
 wire \top_I.branch[21].l_um_ena[9] ;
 wire \top_I.branch[21].l_um_iw[0] ;
 wire \top_I.branch[21].l_um_iw[100] ;
 wire \top_I.branch[21].l_um_iw[101] ;
 wire \top_I.branch[21].l_um_iw[102] ;
 wire \top_I.branch[21].l_um_iw[103] ;
 wire \top_I.branch[21].l_um_iw[104] ;
 wire \top_I.branch[21].l_um_iw[105] ;
 wire \top_I.branch[21].l_um_iw[106] ;
 wire \top_I.branch[21].l_um_iw[107] ;
 wire \top_I.branch[21].l_um_iw[108] ;
 wire \top_I.branch[21].l_um_iw[109] ;
 wire \top_I.branch[21].l_um_iw[10] ;
 wire \top_I.branch[21].l_um_iw[110] ;
 wire \top_I.branch[21].l_um_iw[111] ;
 wire \top_I.branch[21].l_um_iw[112] ;
 wire \top_I.branch[21].l_um_iw[113] ;
 wire \top_I.branch[21].l_um_iw[114] ;
 wire \top_I.branch[21].l_um_iw[115] ;
 wire \top_I.branch[21].l_um_iw[116] ;
 wire \top_I.branch[21].l_um_iw[117] ;
 wire \top_I.branch[21].l_um_iw[118] ;
 wire \top_I.branch[21].l_um_iw[119] ;
 wire \top_I.branch[21].l_um_iw[11] ;
 wire \top_I.branch[21].l_um_iw[120] ;
 wire \top_I.branch[21].l_um_iw[121] ;
 wire \top_I.branch[21].l_um_iw[122] ;
 wire \top_I.branch[21].l_um_iw[123] ;
 wire \top_I.branch[21].l_um_iw[124] ;
 wire \top_I.branch[21].l_um_iw[125] ;
 wire \top_I.branch[21].l_um_iw[126] ;
 wire \top_I.branch[21].l_um_iw[127] ;
 wire \top_I.branch[21].l_um_iw[128] ;
 wire \top_I.branch[21].l_um_iw[129] ;
 wire \top_I.branch[21].l_um_iw[12] ;
 wire \top_I.branch[21].l_um_iw[130] ;
 wire \top_I.branch[21].l_um_iw[131] ;
 wire \top_I.branch[21].l_um_iw[132] ;
 wire \top_I.branch[21].l_um_iw[133] ;
 wire \top_I.branch[21].l_um_iw[134] ;
 wire \top_I.branch[21].l_um_iw[135] ;
 wire \top_I.branch[21].l_um_iw[136] ;
 wire \top_I.branch[21].l_um_iw[137] ;
 wire \top_I.branch[21].l_um_iw[138] ;
 wire \top_I.branch[21].l_um_iw[139] ;
 wire \top_I.branch[21].l_um_iw[13] ;
 wire \top_I.branch[21].l_um_iw[140] ;
 wire \top_I.branch[21].l_um_iw[141] ;
 wire \top_I.branch[21].l_um_iw[142] ;
 wire \top_I.branch[21].l_um_iw[143] ;
 wire \top_I.branch[21].l_um_iw[144] ;
 wire \top_I.branch[21].l_um_iw[145] ;
 wire \top_I.branch[21].l_um_iw[146] ;
 wire \top_I.branch[21].l_um_iw[147] ;
 wire \top_I.branch[21].l_um_iw[148] ;
 wire \top_I.branch[21].l_um_iw[149] ;
 wire \top_I.branch[21].l_um_iw[14] ;
 wire \top_I.branch[21].l_um_iw[150] ;
 wire \top_I.branch[21].l_um_iw[151] ;
 wire \top_I.branch[21].l_um_iw[152] ;
 wire \top_I.branch[21].l_um_iw[153] ;
 wire \top_I.branch[21].l_um_iw[154] ;
 wire \top_I.branch[21].l_um_iw[155] ;
 wire \top_I.branch[21].l_um_iw[156] ;
 wire \top_I.branch[21].l_um_iw[157] ;
 wire \top_I.branch[21].l_um_iw[158] ;
 wire \top_I.branch[21].l_um_iw[159] ;
 wire \top_I.branch[21].l_um_iw[15] ;
 wire \top_I.branch[21].l_um_iw[160] ;
 wire \top_I.branch[21].l_um_iw[161] ;
 wire \top_I.branch[21].l_um_iw[162] ;
 wire \top_I.branch[21].l_um_iw[163] ;
 wire \top_I.branch[21].l_um_iw[164] ;
 wire \top_I.branch[21].l_um_iw[165] ;
 wire \top_I.branch[21].l_um_iw[166] ;
 wire \top_I.branch[21].l_um_iw[167] ;
 wire \top_I.branch[21].l_um_iw[168] ;
 wire \top_I.branch[21].l_um_iw[169] ;
 wire \top_I.branch[21].l_um_iw[16] ;
 wire \top_I.branch[21].l_um_iw[170] ;
 wire \top_I.branch[21].l_um_iw[171] ;
 wire \top_I.branch[21].l_um_iw[172] ;
 wire \top_I.branch[21].l_um_iw[173] ;
 wire \top_I.branch[21].l_um_iw[174] ;
 wire \top_I.branch[21].l_um_iw[175] ;
 wire \top_I.branch[21].l_um_iw[176] ;
 wire \top_I.branch[21].l_um_iw[177] ;
 wire \top_I.branch[21].l_um_iw[178] ;
 wire \top_I.branch[21].l_um_iw[179] ;
 wire \top_I.branch[21].l_um_iw[17] ;
 wire \top_I.branch[21].l_um_iw[180] ;
 wire \top_I.branch[21].l_um_iw[181] ;
 wire \top_I.branch[21].l_um_iw[182] ;
 wire \top_I.branch[21].l_um_iw[183] ;
 wire \top_I.branch[21].l_um_iw[184] ;
 wire \top_I.branch[21].l_um_iw[185] ;
 wire \top_I.branch[21].l_um_iw[186] ;
 wire \top_I.branch[21].l_um_iw[187] ;
 wire \top_I.branch[21].l_um_iw[188] ;
 wire \top_I.branch[21].l_um_iw[189] ;
 wire \top_I.branch[21].l_um_iw[18] ;
 wire \top_I.branch[21].l_um_iw[190] ;
 wire \top_I.branch[21].l_um_iw[191] ;
 wire \top_I.branch[21].l_um_iw[192] ;
 wire \top_I.branch[21].l_um_iw[193] ;
 wire \top_I.branch[21].l_um_iw[194] ;
 wire \top_I.branch[21].l_um_iw[195] ;
 wire \top_I.branch[21].l_um_iw[196] ;
 wire \top_I.branch[21].l_um_iw[197] ;
 wire \top_I.branch[21].l_um_iw[198] ;
 wire \top_I.branch[21].l_um_iw[199] ;
 wire \top_I.branch[21].l_um_iw[19] ;
 wire \top_I.branch[21].l_um_iw[1] ;
 wire \top_I.branch[21].l_um_iw[200] ;
 wire \top_I.branch[21].l_um_iw[201] ;
 wire \top_I.branch[21].l_um_iw[202] ;
 wire \top_I.branch[21].l_um_iw[203] ;
 wire \top_I.branch[21].l_um_iw[204] ;
 wire \top_I.branch[21].l_um_iw[205] ;
 wire \top_I.branch[21].l_um_iw[206] ;
 wire \top_I.branch[21].l_um_iw[207] ;
 wire \top_I.branch[21].l_um_iw[208] ;
 wire \top_I.branch[21].l_um_iw[209] ;
 wire \top_I.branch[21].l_um_iw[20] ;
 wire \top_I.branch[21].l_um_iw[210] ;
 wire \top_I.branch[21].l_um_iw[211] ;
 wire \top_I.branch[21].l_um_iw[212] ;
 wire \top_I.branch[21].l_um_iw[213] ;
 wire \top_I.branch[21].l_um_iw[214] ;
 wire \top_I.branch[21].l_um_iw[215] ;
 wire \top_I.branch[21].l_um_iw[216] ;
 wire \top_I.branch[21].l_um_iw[217] ;
 wire \top_I.branch[21].l_um_iw[218] ;
 wire \top_I.branch[21].l_um_iw[219] ;
 wire \top_I.branch[21].l_um_iw[21] ;
 wire \top_I.branch[21].l_um_iw[220] ;
 wire \top_I.branch[21].l_um_iw[221] ;
 wire \top_I.branch[21].l_um_iw[222] ;
 wire \top_I.branch[21].l_um_iw[223] ;
 wire \top_I.branch[21].l_um_iw[224] ;
 wire \top_I.branch[21].l_um_iw[225] ;
 wire \top_I.branch[21].l_um_iw[226] ;
 wire \top_I.branch[21].l_um_iw[227] ;
 wire \top_I.branch[21].l_um_iw[228] ;
 wire \top_I.branch[21].l_um_iw[229] ;
 wire \top_I.branch[21].l_um_iw[22] ;
 wire \top_I.branch[21].l_um_iw[230] ;
 wire \top_I.branch[21].l_um_iw[231] ;
 wire \top_I.branch[21].l_um_iw[232] ;
 wire \top_I.branch[21].l_um_iw[233] ;
 wire \top_I.branch[21].l_um_iw[234] ;
 wire \top_I.branch[21].l_um_iw[235] ;
 wire \top_I.branch[21].l_um_iw[236] ;
 wire \top_I.branch[21].l_um_iw[237] ;
 wire \top_I.branch[21].l_um_iw[238] ;
 wire \top_I.branch[21].l_um_iw[239] ;
 wire \top_I.branch[21].l_um_iw[23] ;
 wire \top_I.branch[21].l_um_iw[240] ;
 wire \top_I.branch[21].l_um_iw[241] ;
 wire \top_I.branch[21].l_um_iw[242] ;
 wire \top_I.branch[21].l_um_iw[243] ;
 wire \top_I.branch[21].l_um_iw[244] ;
 wire \top_I.branch[21].l_um_iw[245] ;
 wire \top_I.branch[21].l_um_iw[246] ;
 wire \top_I.branch[21].l_um_iw[247] ;
 wire \top_I.branch[21].l_um_iw[248] ;
 wire \top_I.branch[21].l_um_iw[249] ;
 wire \top_I.branch[21].l_um_iw[24] ;
 wire \top_I.branch[21].l_um_iw[250] ;
 wire \top_I.branch[21].l_um_iw[251] ;
 wire \top_I.branch[21].l_um_iw[252] ;
 wire \top_I.branch[21].l_um_iw[253] ;
 wire \top_I.branch[21].l_um_iw[254] ;
 wire \top_I.branch[21].l_um_iw[255] ;
 wire \top_I.branch[21].l_um_iw[256] ;
 wire \top_I.branch[21].l_um_iw[257] ;
 wire \top_I.branch[21].l_um_iw[258] ;
 wire \top_I.branch[21].l_um_iw[259] ;
 wire \top_I.branch[21].l_um_iw[25] ;
 wire \top_I.branch[21].l_um_iw[260] ;
 wire \top_I.branch[21].l_um_iw[261] ;
 wire \top_I.branch[21].l_um_iw[262] ;
 wire \top_I.branch[21].l_um_iw[263] ;
 wire \top_I.branch[21].l_um_iw[264] ;
 wire \top_I.branch[21].l_um_iw[265] ;
 wire \top_I.branch[21].l_um_iw[266] ;
 wire \top_I.branch[21].l_um_iw[267] ;
 wire \top_I.branch[21].l_um_iw[268] ;
 wire \top_I.branch[21].l_um_iw[269] ;
 wire \top_I.branch[21].l_um_iw[26] ;
 wire \top_I.branch[21].l_um_iw[270] ;
 wire \top_I.branch[21].l_um_iw[271] ;
 wire \top_I.branch[21].l_um_iw[272] ;
 wire \top_I.branch[21].l_um_iw[273] ;
 wire \top_I.branch[21].l_um_iw[274] ;
 wire \top_I.branch[21].l_um_iw[275] ;
 wire \top_I.branch[21].l_um_iw[276] ;
 wire \top_I.branch[21].l_um_iw[277] ;
 wire \top_I.branch[21].l_um_iw[278] ;
 wire \top_I.branch[21].l_um_iw[279] ;
 wire \top_I.branch[21].l_um_iw[27] ;
 wire \top_I.branch[21].l_um_iw[280] ;
 wire \top_I.branch[21].l_um_iw[281] ;
 wire \top_I.branch[21].l_um_iw[282] ;
 wire \top_I.branch[21].l_um_iw[283] ;
 wire \top_I.branch[21].l_um_iw[284] ;
 wire \top_I.branch[21].l_um_iw[285] ;
 wire \top_I.branch[21].l_um_iw[286] ;
 wire \top_I.branch[21].l_um_iw[287] ;
 wire \top_I.branch[21].l_um_iw[28] ;
 wire \top_I.branch[21].l_um_iw[29] ;
 wire \top_I.branch[21].l_um_iw[2] ;
 wire \top_I.branch[21].l_um_iw[30] ;
 wire \top_I.branch[21].l_um_iw[31] ;
 wire \top_I.branch[21].l_um_iw[32] ;
 wire \top_I.branch[21].l_um_iw[33] ;
 wire \top_I.branch[21].l_um_iw[34] ;
 wire \top_I.branch[21].l_um_iw[35] ;
 wire \top_I.branch[21].l_um_iw[36] ;
 wire \top_I.branch[21].l_um_iw[37] ;
 wire \top_I.branch[21].l_um_iw[38] ;
 wire \top_I.branch[21].l_um_iw[39] ;
 wire \top_I.branch[21].l_um_iw[3] ;
 wire \top_I.branch[21].l_um_iw[40] ;
 wire \top_I.branch[21].l_um_iw[41] ;
 wire \top_I.branch[21].l_um_iw[42] ;
 wire \top_I.branch[21].l_um_iw[43] ;
 wire \top_I.branch[21].l_um_iw[44] ;
 wire \top_I.branch[21].l_um_iw[45] ;
 wire \top_I.branch[21].l_um_iw[46] ;
 wire \top_I.branch[21].l_um_iw[47] ;
 wire \top_I.branch[21].l_um_iw[48] ;
 wire \top_I.branch[21].l_um_iw[49] ;
 wire \top_I.branch[21].l_um_iw[4] ;
 wire \top_I.branch[21].l_um_iw[50] ;
 wire \top_I.branch[21].l_um_iw[51] ;
 wire \top_I.branch[21].l_um_iw[52] ;
 wire \top_I.branch[21].l_um_iw[53] ;
 wire \top_I.branch[21].l_um_iw[54] ;
 wire \top_I.branch[21].l_um_iw[55] ;
 wire \top_I.branch[21].l_um_iw[56] ;
 wire \top_I.branch[21].l_um_iw[57] ;
 wire \top_I.branch[21].l_um_iw[58] ;
 wire \top_I.branch[21].l_um_iw[59] ;
 wire \top_I.branch[21].l_um_iw[5] ;
 wire \top_I.branch[21].l_um_iw[60] ;
 wire \top_I.branch[21].l_um_iw[61] ;
 wire \top_I.branch[21].l_um_iw[62] ;
 wire \top_I.branch[21].l_um_iw[63] ;
 wire \top_I.branch[21].l_um_iw[64] ;
 wire \top_I.branch[21].l_um_iw[65] ;
 wire \top_I.branch[21].l_um_iw[66] ;
 wire \top_I.branch[21].l_um_iw[67] ;
 wire \top_I.branch[21].l_um_iw[68] ;
 wire \top_I.branch[21].l_um_iw[69] ;
 wire \top_I.branch[21].l_um_iw[6] ;
 wire \top_I.branch[21].l_um_iw[70] ;
 wire \top_I.branch[21].l_um_iw[71] ;
 wire \top_I.branch[21].l_um_iw[72] ;
 wire \top_I.branch[21].l_um_iw[73] ;
 wire \top_I.branch[21].l_um_iw[74] ;
 wire \top_I.branch[21].l_um_iw[75] ;
 wire \top_I.branch[21].l_um_iw[76] ;
 wire \top_I.branch[21].l_um_iw[77] ;
 wire \top_I.branch[21].l_um_iw[78] ;
 wire \top_I.branch[21].l_um_iw[79] ;
 wire \top_I.branch[21].l_um_iw[7] ;
 wire \top_I.branch[21].l_um_iw[80] ;
 wire \top_I.branch[21].l_um_iw[81] ;
 wire \top_I.branch[21].l_um_iw[82] ;
 wire \top_I.branch[21].l_um_iw[83] ;
 wire \top_I.branch[21].l_um_iw[84] ;
 wire \top_I.branch[21].l_um_iw[85] ;
 wire \top_I.branch[21].l_um_iw[86] ;
 wire \top_I.branch[21].l_um_iw[87] ;
 wire \top_I.branch[21].l_um_iw[88] ;
 wire \top_I.branch[21].l_um_iw[89] ;
 wire \top_I.branch[21].l_um_iw[8] ;
 wire \top_I.branch[21].l_um_iw[90] ;
 wire \top_I.branch[21].l_um_iw[91] ;
 wire \top_I.branch[21].l_um_iw[92] ;
 wire \top_I.branch[21].l_um_iw[93] ;
 wire \top_I.branch[21].l_um_iw[94] ;
 wire \top_I.branch[21].l_um_iw[95] ;
 wire \top_I.branch[21].l_um_iw[96] ;
 wire \top_I.branch[21].l_um_iw[97] ;
 wire \top_I.branch[21].l_um_iw[98] ;
 wire \top_I.branch[21].l_um_iw[99] ;
 wire \top_I.branch[21].l_um_iw[9] ;
 wire \top_I.branch[21].l_um_k_zero[0] ;
 wire \top_I.branch[21].l_um_k_zero[10] ;
 wire \top_I.branch[21].l_um_k_zero[11] ;
 wire \top_I.branch[21].l_um_k_zero[12] ;
 wire \top_I.branch[21].l_um_k_zero[13] ;
 wire \top_I.branch[21].l_um_k_zero[14] ;
 wire \top_I.branch[21].l_um_k_zero[15] ;
 wire \top_I.branch[21].l_um_k_zero[1] ;
 wire \top_I.branch[21].l_um_k_zero[2] ;
 wire \top_I.branch[21].l_um_k_zero[3] ;
 wire \top_I.branch[21].l_um_k_zero[4] ;
 wire \top_I.branch[21].l_um_k_zero[5] ;
 wire \top_I.branch[21].l_um_k_zero[6] ;
 wire \top_I.branch[21].l_um_k_zero[7] ;
 wire \top_I.branch[21].l_um_k_zero[8] ;
 wire \top_I.branch[21].l_um_k_zero[9] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[22].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[22].l_k_one ;
 wire \top_I.branch[22].l_k_zero ;
 wire \top_I.branch[22].l_um_ena[0] ;
 wire \top_I.branch[22].l_um_ena[10] ;
 wire \top_I.branch[22].l_um_ena[11] ;
 wire \top_I.branch[22].l_um_ena[12] ;
 wire \top_I.branch[22].l_um_ena[13] ;
 wire \top_I.branch[22].l_um_ena[14] ;
 wire \top_I.branch[22].l_um_ena[15] ;
 wire \top_I.branch[22].l_um_ena[1] ;
 wire \top_I.branch[22].l_um_ena[2] ;
 wire \top_I.branch[22].l_um_ena[3] ;
 wire \top_I.branch[22].l_um_ena[4] ;
 wire \top_I.branch[22].l_um_ena[5] ;
 wire \top_I.branch[22].l_um_ena[6] ;
 wire \top_I.branch[22].l_um_ena[7] ;
 wire \top_I.branch[22].l_um_ena[8] ;
 wire \top_I.branch[22].l_um_ena[9] ;
 wire \top_I.branch[22].l_um_iw[0] ;
 wire \top_I.branch[22].l_um_iw[100] ;
 wire \top_I.branch[22].l_um_iw[101] ;
 wire \top_I.branch[22].l_um_iw[102] ;
 wire \top_I.branch[22].l_um_iw[103] ;
 wire \top_I.branch[22].l_um_iw[104] ;
 wire \top_I.branch[22].l_um_iw[105] ;
 wire \top_I.branch[22].l_um_iw[106] ;
 wire \top_I.branch[22].l_um_iw[107] ;
 wire \top_I.branch[22].l_um_iw[108] ;
 wire \top_I.branch[22].l_um_iw[109] ;
 wire \top_I.branch[22].l_um_iw[10] ;
 wire \top_I.branch[22].l_um_iw[110] ;
 wire \top_I.branch[22].l_um_iw[111] ;
 wire \top_I.branch[22].l_um_iw[112] ;
 wire \top_I.branch[22].l_um_iw[113] ;
 wire \top_I.branch[22].l_um_iw[114] ;
 wire \top_I.branch[22].l_um_iw[115] ;
 wire \top_I.branch[22].l_um_iw[116] ;
 wire \top_I.branch[22].l_um_iw[117] ;
 wire \top_I.branch[22].l_um_iw[118] ;
 wire \top_I.branch[22].l_um_iw[119] ;
 wire \top_I.branch[22].l_um_iw[11] ;
 wire \top_I.branch[22].l_um_iw[120] ;
 wire \top_I.branch[22].l_um_iw[121] ;
 wire \top_I.branch[22].l_um_iw[122] ;
 wire \top_I.branch[22].l_um_iw[123] ;
 wire \top_I.branch[22].l_um_iw[124] ;
 wire \top_I.branch[22].l_um_iw[125] ;
 wire \top_I.branch[22].l_um_iw[126] ;
 wire \top_I.branch[22].l_um_iw[127] ;
 wire \top_I.branch[22].l_um_iw[128] ;
 wire \top_I.branch[22].l_um_iw[129] ;
 wire \top_I.branch[22].l_um_iw[12] ;
 wire \top_I.branch[22].l_um_iw[130] ;
 wire \top_I.branch[22].l_um_iw[131] ;
 wire \top_I.branch[22].l_um_iw[132] ;
 wire \top_I.branch[22].l_um_iw[133] ;
 wire \top_I.branch[22].l_um_iw[134] ;
 wire \top_I.branch[22].l_um_iw[135] ;
 wire \top_I.branch[22].l_um_iw[136] ;
 wire \top_I.branch[22].l_um_iw[137] ;
 wire \top_I.branch[22].l_um_iw[138] ;
 wire \top_I.branch[22].l_um_iw[139] ;
 wire \top_I.branch[22].l_um_iw[13] ;
 wire \top_I.branch[22].l_um_iw[140] ;
 wire \top_I.branch[22].l_um_iw[141] ;
 wire \top_I.branch[22].l_um_iw[142] ;
 wire \top_I.branch[22].l_um_iw[143] ;
 wire \top_I.branch[22].l_um_iw[144] ;
 wire \top_I.branch[22].l_um_iw[145] ;
 wire \top_I.branch[22].l_um_iw[146] ;
 wire \top_I.branch[22].l_um_iw[147] ;
 wire \top_I.branch[22].l_um_iw[148] ;
 wire \top_I.branch[22].l_um_iw[149] ;
 wire \top_I.branch[22].l_um_iw[14] ;
 wire \top_I.branch[22].l_um_iw[150] ;
 wire \top_I.branch[22].l_um_iw[151] ;
 wire \top_I.branch[22].l_um_iw[152] ;
 wire \top_I.branch[22].l_um_iw[153] ;
 wire \top_I.branch[22].l_um_iw[154] ;
 wire \top_I.branch[22].l_um_iw[155] ;
 wire \top_I.branch[22].l_um_iw[156] ;
 wire \top_I.branch[22].l_um_iw[157] ;
 wire \top_I.branch[22].l_um_iw[158] ;
 wire \top_I.branch[22].l_um_iw[159] ;
 wire \top_I.branch[22].l_um_iw[15] ;
 wire \top_I.branch[22].l_um_iw[160] ;
 wire \top_I.branch[22].l_um_iw[161] ;
 wire \top_I.branch[22].l_um_iw[162] ;
 wire \top_I.branch[22].l_um_iw[163] ;
 wire \top_I.branch[22].l_um_iw[164] ;
 wire \top_I.branch[22].l_um_iw[165] ;
 wire \top_I.branch[22].l_um_iw[166] ;
 wire \top_I.branch[22].l_um_iw[167] ;
 wire \top_I.branch[22].l_um_iw[168] ;
 wire \top_I.branch[22].l_um_iw[169] ;
 wire \top_I.branch[22].l_um_iw[16] ;
 wire \top_I.branch[22].l_um_iw[170] ;
 wire \top_I.branch[22].l_um_iw[171] ;
 wire \top_I.branch[22].l_um_iw[172] ;
 wire \top_I.branch[22].l_um_iw[173] ;
 wire \top_I.branch[22].l_um_iw[174] ;
 wire \top_I.branch[22].l_um_iw[175] ;
 wire \top_I.branch[22].l_um_iw[176] ;
 wire \top_I.branch[22].l_um_iw[177] ;
 wire \top_I.branch[22].l_um_iw[178] ;
 wire \top_I.branch[22].l_um_iw[179] ;
 wire \top_I.branch[22].l_um_iw[17] ;
 wire \top_I.branch[22].l_um_iw[180] ;
 wire \top_I.branch[22].l_um_iw[181] ;
 wire \top_I.branch[22].l_um_iw[182] ;
 wire \top_I.branch[22].l_um_iw[183] ;
 wire \top_I.branch[22].l_um_iw[184] ;
 wire \top_I.branch[22].l_um_iw[185] ;
 wire \top_I.branch[22].l_um_iw[186] ;
 wire \top_I.branch[22].l_um_iw[187] ;
 wire \top_I.branch[22].l_um_iw[188] ;
 wire \top_I.branch[22].l_um_iw[189] ;
 wire \top_I.branch[22].l_um_iw[18] ;
 wire \top_I.branch[22].l_um_iw[190] ;
 wire \top_I.branch[22].l_um_iw[191] ;
 wire \top_I.branch[22].l_um_iw[192] ;
 wire \top_I.branch[22].l_um_iw[193] ;
 wire \top_I.branch[22].l_um_iw[194] ;
 wire \top_I.branch[22].l_um_iw[195] ;
 wire \top_I.branch[22].l_um_iw[196] ;
 wire \top_I.branch[22].l_um_iw[197] ;
 wire \top_I.branch[22].l_um_iw[198] ;
 wire \top_I.branch[22].l_um_iw[199] ;
 wire \top_I.branch[22].l_um_iw[19] ;
 wire \top_I.branch[22].l_um_iw[1] ;
 wire \top_I.branch[22].l_um_iw[200] ;
 wire \top_I.branch[22].l_um_iw[201] ;
 wire \top_I.branch[22].l_um_iw[202] ;
 wire \top_I.branch[22].l_um_iw[203] ;
 wire \top_I.branch[22].l_um_iw[204] ;
 wire \top_I.branch[22].l_um_iw[205] ;
 wire \top_I.branch[22].l_um_iw[206] ;
 wire \top_I.branch[22].l_um_iw[207] ;
 wire \top_I.branch[22].l_um_iw[208] ;
 wire \top_I.branch[22].l_um_iw[209] ;
 wire \top_I.branch[22].l_um_iw[20] ;
 wire \top_I.branch[22].l_um_iw[210] ;
 wire \top_I.branch[22].l_um_iw[211] ;
 wire \top_I.branch[22].l_um_iw[212] ;
 wire \top_I.branch[22].l_um_iw[213] ;
 wire \top_I.branch[22].l_um_iw[214] ;
 wire \top_I.branch[22].l_um_iw[215] ;
 wire \top_I.branch[22].l_um_iw[216] ;
 wire \top_I.branch[22].l_um_iw[217] ;
 wire \top_I.branch[22].l_um_iw[218] ;
 wire \top_I.branch[22].l_um_iw[219] ;
 wire \top_I.branch[22].l_um_iw[21] ;
 wire \top_I.branch[22].l_um_iw[220] ;
 wire \top_I.branch[22].l_um_iw[221] ;
 wire \top_I.branch[22].l_um_iw[222] ;
 wire \top_I.branch[22].l_um_iw[223] ;
 wire \top_I.branch[22].l_um_iw[224] ;
 wire \top_I.branch[22].l_um_iw[225] ;
 wire \top_I.branch[22].l_um_iw[226] ;
 wire \top_I.branch[22].l_um_iw[227] ;
 wire \top_I.branch[22].l_um_iw[228] ;
 wire \top_I.branch[22].l_um_iw[229] ;
 wire \top_I.branch[22].l_um_iw[22] ;
 wire \top_I.branch[22].l_um_iw[230] ;
 wire \top_I.branch[22].l_um_iw[231] ;
 wire \top_I.branch[22].l_um_iw[232] ;
 wire \top_I.branch[22].l_um_iw[233] ;
 wire \top_I.branch[22].l_um_iw[234] ;
 wire \top_I.branch[22].l_um_iw[235] ;
 wire \top_I.branch[22].l_um_iw[236] ;
 wire \top_I.branch[22].l_um_iw[237] ;
 wire \top_I.branch[22].l_um_iw[238] ;
 wire \top_I.branch[22].l_um_iw[239] ;
 wire \top_I.branch[22].l_um_iw[23] ;
 wire \top_I.branch[22].l_um_iw[240] ;
 wire \top_I.branch[22].l_um_iw[241] ;
 wire \top_I.branch[22].l_um_iw[242] ;
 wire \top_I.branch[22].l_um_iw[243] ;
 wire \top_I.branch[22].l_um_iw[244] ;
 wire \top_I.branch[22].l_um_iw[245] ;
 wire \top_I.branch[22].l_um_iw[246] ;
 wire \top_I.branch[22].l_um_iw[247] ;
 wire \top_I.branch[22].l_um_iw[248] ;
 wire \top_I.branch[22].l_um_iw[249] ;
 wire \top_I.branch[22].l_um_iw[24] ;
 wire \top_I.branch[22].l_um_iw[250] ;
 wire \top_I.branch[22].l_um_iw[251] ;
 wire \top_I.branch[22].l_um_iw[252] ;
 wire \top_I.branch[22].l_um_iw[253] ;
 wire \top_I.branch[22].l_um_iw[254] ;
 wire \top_I.branch[22].l_um_iw[255] ;
 wire \top_I.branch[22].l_um_iw[256] ;
 wire \top_I.branch[22].l_um_iw[257] ;
 wire \top_I.branch[22].l_um_iw[258] ;
 wire \top_I.branch[22].l_um_iw[259] ;
 wire \top_I.branch[22].l_um_iw[25] ;
 wire \top_I.branch[22].l_um_iw[260] ;
 wire \top_I.branch[22].l_um_iw[261] ;
 wire \top_I.branch[22].l_um_iw[262] ;
 wire \top_I.branch[22].l_um_iw[263] ;
 wire \top_I.branch[22].l_um_iw[264] ;
 wire \top_I.branch[22].l_um_iw[265] ;
 wire \top_I.branch[22].l_um_iw[266] ;
 wire \top_I.branch[22].l_um_iw[267] ;
 wire \top_I.branch[22].l_um_iw[268] ;
 wire \top_I.branch[22].l_um_iw[269] ;
 wire \top_I.branch[22].l_um_iw[26] ;
 wire \top_I.branch[22].l_um_iw[270] ;
 wire \top_I.branch[22].l_um_iw[271] ;
 wire \top_I.branch[22].l_um_iw[272] ;
 wire \top_I.branch[22].l_um_iw[273] ;
 wire \top_I.branch[22].l_um_iw[274] ;
 wire \top_I.branch[22].l_um_iw[275] ;
 wire \top_I.branch[22].l_um_iw[276] ;
 wire \top_I.branch[22].l_um_iw[277] ;
 wire \top_I.branch[22].l_um_iw[278] ;
 wire \top_I.branch[22].l_um_iw[279] ;
 wire \top_I.branch[22].l_um_iw[27] ;
 wire \top_I.branch[22].l_um_iw[280] ;
 wire \top_I.branch[22].l_um_iw[281] ;
 wire \top_I.branch[22].l_um_iw[282] ;
 wire \top_I.branch[22].l_um_iw[283] ;
 wire \top_I.branch[22].l_um_iw[284] ;
 wire \top_I.branch[22].l_um_iw[285] ;
 wire \top_I.branch[22].l_um_iw[286] ;
 wire \top_I.branch[22].l_um_iw[287] ;
 wire \top_I.branch[22].l_um_iw[28] ;
 wire \top_I.branch[22].l_um_iw[29] ;
 wire \top_I.branch[22].l_um_iw[2] ;
 wire \top_I.branch[22].l_um_iw[30] ;
 wire \top_I.branch[22].l_um_iw[31] ;
 wire \top_I.branch[22].l_um_iw[32] ;
 wire \top_I.branch[22].l_um_iw[33] ;
 wire \top_I.branch[22].l_um_iw[34] ;
 wire \top_I.branch[22].l_um_iw[35] ;
 wire \top_I.branch[22].l_um_iw[36] ;
 wire \top_I.branch[22].l_um_iw[37] ;
 wire \top_I.branch[22].l_um_iw[38] ;
 wire \top_I.branch[22].l_um_iw[39] ;
 wire \top_I.branch[22].l_um_iw[3] ;
 wire \top_I.branch[22].l_um_iw[40] ;
 wire \top_I.branch[22].l_um_iw[41] ;
 wire \top_I.branch[22].l_um_iw[42] ;
 wire \top_I.branch[22].l_um_iw[43] ;
 wire \top_I.branch[22].l_um_iw[44] ;
 wire \top_I.branch[22].l_um_iw[45] ;
 wire \top_I.branch[22].l_um_iw[46] ;
 wire \top_I.branch[22].l_um_iw[47] ;
 wire \top_I.branch[22].l_um_iw[48] ;
 wire \top_I.branch[22].l_um_iw[49] ;
 wire \top_I.branch[22].l_um_iw[4] ;
 wire \top_I.branch[22].l_um_iw[50] ;
 wire \top_I.branch[22].l_um_iw[51] ;
 wire \top_I.branch[22].l_um_iw[52] ;
 wire \top_I.branch[22].l_um_iw[53] ;
 wire \top_I.branch[22].l_um_iw[54] ;
 wire \top_I.branch[22].l_um_iw[55] ;
 wire \top_I.branch[22].l_um_iw[56] ;
 wire \top_I.branch[22].l_um_iw[57] ;
 wire \top_I.branch[22].l_um_iw[58] ;
 wire \top_I.branch[22].l_um_iw[59] ;
 wire \top_I.branch[22].l_um_iw[5] ;
 wire \top_I.branch[22].l_um_iw[60] ;
 wire \top_I.branch[22].l_um_iw[61] ;
 wire \top_I.branch[22].l_um_iw[62] ;
 wire \top_I.branch[22].l_um_iw[63] ;
 wire \top_I.branch[22].l_um_iw[64] ;
 wire \top_I.branch[22].l_um_iw[65] ;
 wire \top_I.branch[22].l_um_iw[66] ;
 wire \top_I.branch[22].l_um_iw[67] ;
 wire \top_I.branch[22].l_um_iw[68] ;
 wire \top_I.branch[22].l_um_iw[69] ;
 wire \top_I.branch[22].l_um_iw[6] ;
 wire \top_I.branch[22].l_um_iw[70] ;
 wire \top_I.branch[22].l_um_iw[71] ;
 wire \top_I.branch[22].l_um_iw[72] ;
 wire \top_I.branch[22].l_um_iw[73] ;
 wire \top_I.branch[22].l_um_iw[74] ;
 wire \top_I.branch[22].l_um_iw[75] ;
 wire \top_I.branch[22].l_um_iw[76] ;
 wire \top_I.branch[22].l_um_iw[77] ;
 wire \top_I.branch[22].l_um_iw[78] ;
 wire \top_I.branch[22].l_um_iw[79] ;
 wire \top_I.branch[22].l_um_iw[7] ;
 wire \top_I.branch[22].l_um_iw[80] ;
 wire \top_I.branch[22].l_um_iw[81] ;
 wire \top_I.branch[22].l_um_iw[82] ;
 wire \top_I.branch[22].l_um_iw[83] ;
 wire \top_I.branch[22].l_um_iw[84] ;
 wire \top_I.branch[22].l_um_iw[85] ;
 wire \top_I.branch[22].l_um_iw[86] ;
 wire \top_I.branch[22].l_um_iw[87] ;
 wire \top_I.branch[22].l_um_iw[88] ;
 wire \top_I.branch[22].l_um_iw[89] ;
 wire \top_I.branch[22].l_um_iw[8] ;
 wire \top_I.branch[22].l_um_iw[90] ;
 wire \top_I.branch[22].l_um_iw[91] ;
 wire \top_I.branch[22].l_um_iw[92] ;
 wire \top_I.branch[22].l_um_iw[93] ;
 wire \top_I.branch[22].l_um_iw[94] ;
 wire \top_I.branch[22].l_um_iw[95] ;
 wire \top_I.branch[22].l_um_iw[96] ;
 wire \top_I.branch[22].l_um_iw[97] ;
 wire \top_I.branch[22].l_um_iw[98] ;
 wire \top_I.branch[22].l_um_iw[99] ;
 wire \top_I.branch[22].l_um_iw[9] ;
 wire \top_I.branch[22].l_um_k_zero[0] ;
 wire \top_I.branch[22].l_um_k_zero[10] ;
 wire \top_I.branch[22].l_um_k_zero[11] ;
 wire \top_I.branch[22].l_um_k_zero[12] ;
 wire \top_I.branch[22].l_um_k_zero[13] ;
 wire \top_I.branch[22].l_um_k_zero[14] ;
 wire \top_I.branch[22].l_um_k_zero[15] ;
 wire \top_I.branch[22].l_um_k_zero[1] ;
 wire \top_I.branch[22].l_um_k_zero[2] ;
 wire \top_I.branch[22].l_um_k_zero[3] ;
 wire \top_I.branch[22].l_um_k_zero[4] ;
 wire \top_I.branch[22].l_um_k_zero[5] ;
 wire \top_I.branch[22].l_um_k_zero[6] ;
 wire \top_I.branch[22].l_um_k_zero[7] ;
 wire \top_I.branch[22].l_um_k_zero[8] ;
 wire \top_I.branch[22].l_um_k_zero[9] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[23].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[23].l_k_one ;
 wire \top_I.branch[23].l_k_zero ;
 wire \top_I.branch[23].l_um_ena[0] ;
 wire \top_I.branch[23].l_um_ena[10] ;
 wire \top_I.branch[23].l_um_ena[11] ;
 wire \top_I.branch[23].l_um_ena[12] ;
 wire \top_I.branch[23].l_um_ena[13] ;
 wire \top_I.branch[23].l_um_ena[14] ;
 wire \top_I.branch[23].l_um_ena[15] ;
 wire \top_I.branch[23].l_um_ena[1] ;
 wire \top_I.branch[23].l_um_ena[2] ;
 wire \top_I.branch[23].l_um_ena[3] ;
 wire \top_I.branch[23].l_um_ena[4] ;
 wire \top_I.branch[23].l_um_ena[5] ;
 wire \top_I.branch[23].l_um_ena[6] ;
 wire \top_I.branch[23].l_um_ena[7] ;
 wire \top_I.branch[23].l_um_ena[8] ;
 wire \top_I.branch[23].l_um_ena[9] ;
 wire \top_I.branch[23].l_um_iw[0] ;
 wire \top_I.branch[23].l_um_iw[100] ;
 wire \top_I.branch[23].l_um_iw[101] ;
 wire \top_I.branch[23].l_um_iw[102] ;
 wire \top_I.branch[23].l_um_iw[103] ;
 wire \top_I.branch[23].l_um_iw[104] ;
 wire \top_I.branch[23].l_um_iw[105] ;
 wire \top_I.branch[23].l_um_iw[106] ;
 wire \top_I.branch[23].l_um_iw[107] ;
 wire \top_I.branch[23].l_um_iw[108] ;
 wire \top_I.branch[23].l_um_iw[109] ;
 wire \top_I.branch[23].l_um_iw[10] ;
 wire \top_I.branch[23].l_um_iw[110] ;
 wire \top_I.branch[23].l_um_iw[111] ;
 wire \top_I.branch[23].l_um_iw[112] ;
 wire \top_I.branch[23].l_um_iw[113] ;
 wire \top_I.branch[23].l_um_iw[114] ;
 wire \top_I.branch[23].l_um_iw[115] ;
 wire \top_I.branch[23].l_um_iw[116] ;
 wire \top_I.branch[23].l_um_iw[117] ;
 wire \top_I.branch[23].l_um_iw[118] ;
 wire \top_I.branch[23].l_um_iw[119] ;
 wire \top_I.branch[23].l_um_iw[11] ;
 wire \top_I.branch[23].l_um_iw[120] ;
 wire \top_I.branch[23].l_um_iw[121] ;
 wire \top_I.branch[23].l_um_iw[122] ;
 wire \top_I.branch[23].l_um_iw[123] ;
 wire \top_I.branch[23].l_um_iw[124] ;
 wire \top_I.branch[23].l_um_iw[125] ;
 wire \top_I.branch[23].l_um_iw[126] ;
 wire \top_I.branch[23].l_um_iw[127] ;
 wire \top_I.branch[23].l_um_iw[128] ;
 wire \top_I.branch[23].l_um_iw[129] ;
 wire \top_I.branch[23].l_um_iw[12] ;
 wire \top_I.branch[23].l_um_iw[130] ;
 wire \top_I.branch[23].l_um_iw[131] ;
 wire \top_I.branch[23].l_um_iw[132] ;
 wire \top_I.branch[23].l_um_iw[133] ;
 wire \top_I.branch[23].l_um_iw[134] ;
 wire \top_I.branch[23].l_um_iw[135] ;
 wire \top_I.branch[23].l_um_iw[136] ;
 wire \top_I.branch[23].l_um_iw[137] ;
 wire \top_I.branch[23].l_um_iw[138] ;
 wire \top_I.branch[23].l_um_iw[139] ;
 wire \top_I.branch[23].l_um_iw[13] ;
 wire \top_I.branch[23].l_um_iw[140] ;
 wire \top_I.branch[23].l_um_iw[141] ;
 wire \top_I.branch[23].l_um_iw[142] ;
 wire \top_I.branch[23].l_um_iw[143] ;
 wire \top_I.branch[23].l_um_iw[144] ;
 wire \top_I.branch[23].l_um_iw[145] ;
 wire \top_I.branch[23].l_um_iw[146] ;
 wire \top_I.branch[23].l_um_iw[147] ;
 wire \top_I.branch[23].l_um_iw[148] ;
 wire \top_I.branch[23].l_um_iw[149] ;
 wire \top_I.branch[23].l_um_iw[14] ;
 wire \top_I.branch[23].l_um_iw[150] ;
 wire \top_I.branch[23].l_um_iw[151] ;
 wire \top_I.branch[23].l_um_iw[152] ;
 wire \top_I.branch[23].l_um_iw[153] ;
 wire \top_I.branch[23].l_um_iw[154] ;
 wire \top_I.branch[23].l_um_iw[155] ;
 wire \top_I.branch[23].l_um_iw[156] ;
 wire \top_I.branch[23].l_um_iw[157] ;
 wire \top_I.branch[23].l_um_iw[158] ;
 wire \top_I.branch[23].l_um_iw[159] ;
 wire \top_I.branch[23].l_um_iw[15] ;
 wire \top_I.branch[23].l_um_iw[160] ;
 wire \top_I.branch[23].l_um_iw[161] ;
 wire \top_I.branch[23].l_um_iw[162] ;
 wire \top_I.branch[23].l_um_iw[163] ;
 wire \top_I.branch[23].l_um_iw[164] ;
 wire \top_I.branch[23].l_um_iw[165] ;
 wire \top_I.branch[23].l_um_iw[166] ;
 wire \top_I.branch[23].l_um_iw[167] ;
 wire \top_I.branch[23].l_um_iw[168] ;
 wire \top_I.branch[23].l_um_iw[169] ;
 wire \top_I.branch[23].l_um_iw[16] ;
 wire \top_I.branch[23].l_um_iw[170] ;
 wire \top_I.branch[23].l_um_iw[171] ;
 wire \top_I.branch[23].l_um_iw[172] ;
 wire \top_I.branch[23].l_um_iw[173] ;
 wire \top_I.branch[23].l_um_iw[174] ;
 wire \top_I.branch[23].l_um_iw[175] ;
 wire \top_I.branch[23].l_um_iw[176] ;
 wire \top_I.branch[23].l_um_iw[177] ;
 wire \top_I.branch[23].l_um_iw[178] ;
 wire \top_I.branch[23].l_um_iw[179] ;
 wire \top_I.branch[23].l_um_iw[17] ;
 wire \top_I.branch[23].l_um_iw[180] ;
 wire \top_I.branch[23].l_um_iw[181] ;
 wire \top_I.branch[23].l_um_iw[182] ;
 wire \top_I.branch[23].l_um_iw[183] ;
 wire \top_I.branch[23].l_um_iw[184] ;
 wire \top_I.branch[23].l_um_iw[185] ;
 wire \top_I.branch[23].l_um_iw[186] ;
 wire \top_I.branch[23].l_um_iw[187] ;
 wire \top_I.branch[23].l_um_iw[188] ;
 wire \top_I.branch[23].l_um_iw[189] ;
 wire \top_I.branch[23].l_um_iw[18] ;
 wire \top_I.branch[23].l_um_iw[190] ;
 wire \top_I.branch[23].l_um_iw[191] ;
 wire \top_I.branch[23].l_um_iw[192] ;
 wire \top_I.branch[23].l_um_iw[193] ;
 wire \top_I.branch[23].l_um_iw[194] ;
 wire \top_I.branch[23].l_um_iw[195] ;
 wire \top_I.branch[23].l_um_iw[196] ;
 wire \top_I.branch[23].l_um_iw[197] ;
 wire \top_I.branch[23].l_um_iw[198] ;
 wire \top_I.branch[23].l_um_iw[199] ;
 wire \top_I.branch[23].l_um_iw[19] ;
 wire \top_I.branch[23].l_um_iw[1] ;
 wire \top_I.branch[23].l_um_iw[200] ;
 wire \top_I.branch[23].l_um_iw[201] ;
 wire \top_I.branch[23].l_um_iw[202] ;
 wire \top_I.branch[23].l_um_iw[203] ;
 wire \top_I.branch[23].l_um_iw[204] ;
 wire \top_I.branch[23].l_um_iw[205] ;
 wire \top_I.branch[23].l_um_iw[206] ;
 wire \top_I.branch[23].l_um_iw[207] ;
 wire \top_I.branch[23].l_um_iw[208] ;
 wire \top_I.branch[23].l_um_iw[209] ;
 wire \top_I.branch[23].l_um_iw[20] ;
 wire \top_I.branch[23].l_um_iw[210] ;
 wire \top_I.branch[23].l_um_iw[211] ;
 wire \top_I.branch[23].l_um_iw[212] ;
 wire \top_I.branch[23].l_um_iw[213] ;
 wire \top_I.branch[23].l_um_iw[214] ;
 wire \top_I.branch[23].l_um_iw[215] ;
 wire \top_I.branch[23].l_um_iw[216] ;
 wire \top_I.branch[23].l_um_iw[217] ;
 wire \top_I.branch[23].l_um_iw[218] ;
 wire \top_I.branch[23].l_um_iw[219] ;
 wire \top_I.branch[23].l_um_iw[21] ;
 wire \top_I.branch[23].l_um_iw[220] ;
 wire \top_I.branch[23].l_um_iw[221] ;
 wire \top_I.branch[23].l_um_iw[222] ;
 wire \top_I.branch[23].l_um_iw[223] ;
 wire \top_I.branch[23].l_um_iw[224] ;
 wire \top_I.branch[23].l_um_iw[225] ;
 wire \top_I.branch[23].l_um_iw[226] ;
 wire \top_I.branch[23].l_um_iw[227] ;
 wire \top_I.branch[23].l_um_iw[228] ;
 wire \top_I.branch[23].l_um_iw[229] ;
 wire \top_I.branch[23].l_um_iw[22] ;
 wire \top_I.branch[23].l_um_iw[230] ;
 wire \top_I.branch[23].l_um_iw[231] ;
 wire \top_I.branch[23].l_um_iw[232] ;
 wire \top_I.branch[23].l_um_iw[233] ;
 wire \top_I.branch[23].l_um_iw[234] ;
 wire \top_I.branch[23].l_um_iw[235] ;
 wire \top_I.branch[23].l_um_iw[236] ;
 wire \top_I.branch[23].l_um_iw[237] ;
 wire \top_I.branch[23].l_um_iw[238] ;
 wire \top_I.branch[23].l_um_iw[239] ;
 wire \top_I.branch[23].l_um_iw[23] ;
 wire \top_I.branch[23].l_um_iw[240] ;
 wire \top_I.branch[23].l_um_iw[241] ;
 wire \top_I.branch[23].l_um_iw[242] ;
 wire \top_I.branch[23].l_um_iw[243] ;
 wire \top_I.branch[23].l_um_iw[244] ;
 wire \top_I.branch[23].l_um_iw[245] ;
 wire \top_I.branch[23].l_um_iw[246] ;
 wire \top_I.branch[23].l_um_iw[247] ;
 wire \top_I.branch[23].l_um_iw[248] ;
 wire \top_I.branch[23].l_um_iw[249] ;
 wire \top_I.branch[23].l_um_iw[24] ;
 wire \top_I.branch[23].l_um_iw[250] ;
 wire \top_I.branch[23].l_um_iw[251] ;
 wire \top_I.branch[23].l_um_iw[252] ;
 wire \top_I.branch[23].l_um_iw[253] ;
 wire \top_I.branch[23].l_um_iw[254] ;
 wire \top_I.branch[23].l_um_iw[255] ;
 wire \top_I.branch[23].l_um_iw[256] ;
 wire \top_I.branch[23].l_um_iw[257] ;
 wire \top_I.branch[23].l_um_iw[258] ;
 wire \top_I.branch[23].l_um_iw[259] ;
 wire \top_I.branch[23].l_um_iw[25] ;
 wire \top_I.branch[23].l_um_iw[260] ;
 wire \top_I.branch[23].l_um_iw[261] ;
 wire \top_I.branch[23].l_um_iw[262] ;
 wire \top_I.branch[23].l_um_iw[263] ;
 wire \top_I.branch[23].l_um_iw[264] ;
 wire \top_I.branch[23].l_um_iw[265] ;
 wire \top_I.branch[23].l_um_iw[266] ;
 wire \top_I.branch[23].l_um_iw[267] ;
 wire \top_I.branch[23].l_um_iw[268] ;
 wire \top_I.branch[23].l_um_iw[269] ;
 wire \top_I.branch[23].l_um_iw[26] ;
 wire \top_I.branch[23].l_um_iw[270] ;
 wire \top_I.branch[23].l_um_iw[271] ;
 wire \top_I.branch[23].l_um_iw[272] ;
 wire \top_I.branch[23].l_um_iw[273] ;
 wire \top_I.branch[23].l_um_iw[274] ;
 wire \top_I.branch[23].l_um_iw[275] ;
 wire \top_I.branch[23].l_um_iw[276] ;
 wire \top_I.branch[23].l_um_iw[277] ;
 wire \top_I.branch[23].l_um_iw[278] ;
 wire \top_I.branch[23].l_um_iw[279] ;
 wire \top_I.branch[23].l_um_iw[27] ;
 wire \top_I.branch[23].l_um_iw[280] ;
 wire \top_I.branch[23].l_um_iw[281] ;
 wire \top_I.branch[23].l_um_iw[282] ;
 wire \top_I.branch[23].l_um_iw[283] ;
 wire \top_I.branch[23].l_um_iw[284] ;
 wire \top_I.branch[23].l_um_iw[285] ;
 wire \top_I.branch[23].l_um_iw[286] ;
 wire \top_I.branch[23].l_um_iw[287] ;
 wire \top_I.branch[23].l_um_iw[28] ;
 wire \top_I.branch[23].l_um_iw[29] ;
 wire \top_I.branch[23].l_um_iw[2] ;
 wire \top_I.branch[23].l_um_iw[30] ;
 wire \top_I.branch[23].l_um_iw[31] ;
 wire \top_I.branch[23].l_um_iw[32] ;
 wire \top_I.branch[23].l_um_iw[33] ;
 wire \top_I.branch[23].l_um_iw[34] ;
 wire \top_I.branch[23].l_um_iw[35] ;
 wire \top_I.branch[23].l_um_iw[36] ;
 wire \top_I.branch[23].l_um_iw[37] ;
 wire \top_I.branch[23].l_um_iw[38] ;
 wire \top_I.branch[23].l_um_iw[39] ;
 wire \top_I.branch[23].l_um_iw[3] ;
 wire \top_I.branch[23].l_um_iw[40] ;
 wire \top_I.branch[23].l_um_iw[41] ;
 wire \top_I.branch[23].l_um_iw[42] ;
 wire \top_I.branch[23].l_um_iw[43] ;
 wire \top_I.branch[23].l_um_iw[44] ;
 wire \top_I.branch[23].l_um_iw[45] ;
 wire \top_I.branch[23].l_um_iw[46] ;
 wire \top_I.branch[23].l_um_iw[47] ;
 wire \top_I.branch[23].l_um_iw[48] ;
 wire \top_I.branch[23].l_um_iw[49] ;
 wire \top_I.branch[23].l_um_iw[4] ;
 wire \top_I.branch[23].l_um_iw[50] ;
 wire \top_I.branch[23].l_um_iw[51] ;
 wire \top_I.branch[23].l_um_iw[52] ;
 wire \top_I.branch[23].l_um_iw[53] ;
 wire \top_I.branch[23].l_um_iw[54] ;
 wire \top_I.branch[23].l_um_iw[55] ;
 wire \top_I.branch[23].l_um_iw[56] ;
 wire \top_I.branch[23].l_um_iw[57] ;
 wire \top_I.branch[23].l_um_iw[58] ;
 wire \top_I.branch[23].l_um_iw[59] ;
 wire \top_I.branch[23].l_um_iw[5] ;
 wire \top_I.branch[23].l_um_iw[60] ;
 wire \top_I.branch[23].l_um_iw[61] ;
 wire \top_I.branch[23].l_um_iw[62] ;
 wire \top_I.branch[23].l_um_iw[63] ;
 wire \top_I.branch[23].l_um_iw[64] ;
 wire \top_I.branch[23].l_um_iw[65] ;
 wire \top_I.branch[23].l_um_iw[66] ;
 wire \top_I.branch[23].l_um_iw[67] ;
 wire \top_I.branch[23].l_um_iw[68] ;
 wire \top_I.branch[23].l_um_iw[69] ;
 wire \top_I.branch[23].l_um_iw[6] ;
 wire \top_I.branch[23].l_um_iw[70] ;
 wire \top_I.branch[23].l_um_iw[71] ;
 wire \top_I.branch[23].l_um_iw[72] ;
 wire \top_I.branch[23].l_um_iw[73] ;
 wire \top_I.branch[23].l_um_iw[74] ;
 wire \top_I.branch[23].l_um_iw[75] ;
 wire \top_I.branch[23].l_um_iw[76] ;
 wire \top_I.branch[23].l_um_iw[77] ;
 wire \top_I.branch[23].l_um_iw[78] ;
 wire \top_I.branch[23].l_um_iw[79] ;
 wire \top_I.branch[23].l_um_iw[7] ;
 wire \top_I.branch[23].l_um_iw[80] ;
 wire \top_I.branch[23].l_um_iw[81] ;
 wire \top_I.branch[23].l_um_iw[82] ;
 wire \top_I.branch[23].l_um_iw[83] ;
 wire \top_I.branch[23].l_um_iw[84] ;
 wire \top_I.branch[23].l_um_iw[85] ;
 wire \top_I.branch[23].l_um_iw[86] ;
 wire \top_I.branch[23].l_um_iw[87] ;
 wire \top_I.branch[23].l_um_iw[88] ;
 wire \top_I.branch[23].l_um_iw[89] ;
 wire \top_I.branch[23].l_um_iw[8] ;
 wire \top_I.branch[23].l_um_iw[90] ;
 wire \top_I.branch[23].l_um_iw[91] ;
 wire \top_I.branch[23].l_um_iw[92] ;
 wire \top_I.branch[23].l_um_iw[93] ;
 wire \top_I.branch[23].l_um_iw[94] ;
 wire \top_I.branch[23].l_um_iw[95] ;
 wire \top_I.branch[23].l_um_iw[96] ;
 wire \top_I.branch[23].l_um_iw[97] ;
 wire \top_I.branch[23].l_um_iw[98] ;
 wire \top_I.branch[23].l_um_iw[99] ;
 wire \top_I.branch[23].l_um_iw[9] ;
 wire \top_I.branch[23].l_um_k_zero[0] ;
 wire \top_I.branch[23].l_um_k_zero[10] ;
 wire \top_I.branch[23].l_um_k_zero[11] ;
 wire \top_I.branch[23].l_um_k_zero[12] ;
 wire \top_I.branch[23].l_um_k_zero[13] ;
 wire \top_I.branch[23].l_um_k_zero[14] ;
 wire \top_I.branch[23].l_um_k_zero[15] ;
 wire \top_I.branch[23].l_um_k_zero[1] ;
 wire \top_I.branch[23].l_um_k_zero[2] ;
 wire \top_I.branch[23].l_um_k_zero[3] ;
 wire \top_I.branch[23].l_um_k_zero[4] ;
 wire \top_I.branch[23].l_um_k_zero[5] ;
 wire \top_I.branch[23].l_um_k_zero[6] ;
 wire \top_I.branch[23].l_um_k_zero[7] ;
 wire \top_I.branch[23].l_um_k_zero[8] ;
 wire \top_I.branch[23].l_um_k_zero[9] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[1].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[2].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[3].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[4].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[5].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[0] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[1] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[2] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[3] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[4] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[5] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[6] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_oe[7] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[0] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[1] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[2] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[3] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[4] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[5] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[6] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uio_out[7] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[0] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[1] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[2] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[3] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[4] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[5] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[6] ;
 wire \top_I.branch[2].col_um[6].um_top_I.uo_out[7] ;
 wire \top_I.branch[2].l_k_one ;
 wire \top_I.branch[2].l_k_zero ;
 wire \top_I.branch[2].l_um_ena[0] ;
 wire \top_I.branch[2].l_um_ena[10] ;
 wire \top_I.branch[2].l_um_ena[11] ;
 wire \top_I.branch[2].l_um_ena[12] ;
 wire \top_I.branch[2].l_um_ena[13] ;
 wire \top_I.branch[2].l_um_ena[14] ;
 wire \top_I.branch[2].l_um_ena[15] ;
 wire \top_I.branch[2].l_um_ena[1] ;
 wire \top_I.branch[2].l_um_ena[2] ;
 wire \top_I.branch[2].l_um_ena[3] ;
 wire \top_I.branch[2].l_um_ena[4] ;
 wire \top_I.branch[2].l_um_ena[5] ;
 wire \top_I.branch[2].l_um_ena[6] ;
 wire \top_I.branch[2].l_um_ena[7] ;
 wire \top_I.branch[2].l_um_ena[8] ;
 wire \top_I.branch[2].l_um_ena[9] ;
 wire \top_I.branch[2].l_um_iw[0] ;
 wire \top_I.branch[2].l_um_iw[100] ;
 wire \top_I.branch[2].l_um_iw[101] ;
 wire \top_I.branch[2].l_um_iw[102] ;
 wire \top_I.branch[2].l_um_iw[103] ;
 wire \top_I.branch[2].l_um_iw[104] ;
 wire \top_I.branch[2].l_um_iw[105] ;
 wire \top_I.branch[2].l_um_iw[106] ;
 wire \top_I.branch[2].l_um_iw[107] ;
 wire \top_I.branch[2].l_um_iw[108] ;
 wire \top_I.branch[2].l_um_iw[109] ;
 wire \top_I.branch[2].l_um_iw[10] ;
 wire \top_I.branch[2].l_um_iw[110] ;
 wire \top_I.branch[2].l_um_iw[111] ;
 wire \top_I.branch[2].l_um_iw[112] ;
 wire \top_I.branch[2].l_um_iw[113] ;
 wire \top_I.branch[2].l_um_iw[114] ;
 wire \top_I.branch[2].l_um_iw[115] ;
 wire \top_I.branch[2].l_um_iw[116] ;
 wire \top_I.branch[2].l_um_iw[117] ;
 wire \top_I.branch[2].l_um_iw[118] ;
 wire \top_I.branch[2].l_um_iw[119] ;
 wire \top_I.branch[2].l_um_iw[11] ;
 wire \top_I.branch[2].l_um_iw[120] ;
 wire \top_I.branch[2].l_um_iw[121] ;
 wire \top_I.branch[2].l_um_iw[122] ;
 wire \top_I.branch[2].l_um_iw[123] ;
 wire \top_I.branch[2].l_um_iw[124] ;
 wire \top_I.branch[2].l_um_iw[125] ;
 wire \top_I.branch[2].l_um_iw[126] ;
 wire \top_I.branch[2].l_um_iw[127] ;
 wire \top_I.branch[2].l_um_iw[128] ;
 wire \top_I.branch[2].l_um_iw[129] ;
 wire \top_I.branch[2].l_um_iw[12] ;
 wire \top_I.branch[2].l_um_iw[130] ;
 wire \top_I.branch[2].l_um_iw[131] ;
 wire \top_I.branch[2].l_um_iw[132] ;
 wire \top_I.branch[2].l_um_iw[133] ;
 wire \top_I.branch[2].l_um_iw[134] ;
 wire \top_I.branch[2].l_um_iw[135] ;
 wire \top_I.branch[2].l_um_iw[136] ;
 wire \top_I.branch[2].l_um_iw[137] ;
 wire \top_I.branch[2].l_um_iw[138] ;
 wire \top_I.branch[2].l_um_iw[139] ;
 wire \top_I.branch[2].l_um_iw[13] ;
 wire \top_I.branch[2].l_um_iw[140] ;
 wire \top_I.branch[2].l_um_iw[141] ;
 wire \top_I.branch[2].l_um_iw[142] ;
 wire \top_I.branch[2].l_um_iw[143] ;
 wire \top_I.branch[2].l_um_iw[144] ;
 wire \top_I.branch[2].l_um_iw[145] ;
 wire \top_I.branch[2].l_um_iw[146] ;
 wire \top_I.branch[2].l_um_iw[147] ;
 wire \top_I.branch[2].l_um_iw[148] ;
 wire \top_I.branch[2].l_um_iw[149] ;
 wire \top_I.branch[2].l_um_iw[14] ;
 wire \top_I.branch[2].l_um_iw[150] ;
 wire \top_I.branch[2].l_um_iw[151] ;
 wire \top_I.branch[2].l_um_iw[152] ;
 wire \top_I.branch[2].l_um_iw[153] ;
 wire \top_I.branch[2].l_um_iw[154] ;
 wire \top_I.branch[2].l_um_iw[155] ;
 wire \top_I.branch[2].l_um_iw[156] ;
 wire \top_I.branch[2].l_um_iw[157] ;
 wire \top_I.branch[2].l_um_iw[158] ;
 wire \top_I.branch[2].l_um_iw[159] ;
 wire \top_I.branch[2].l_um_iw[15] ;
 wire \top_I.branch[2].l_um_iw[160] ;
 wire \top_I.branch[2].l_um_iw[161] ;
 wire \top_I.branch[2].l_um_iw[162] ;
 wire \top_I.branch[2].l_um_iw[163] ;
 wire \top_I.branch[2].l_um_iw[164] ;
 wire \top_I.branch[2].l_um_iw[165] ;
 wire \top_I.branch[2].l_um_iw[166] ;
 wire \top_I.branch[2].l_um_iw[167] ;
 wire \top_I.branch[2].l_um_iw[168] ;
 wire \top_I.branch[2].l_um_iw[169] ;
 wire \top_I.branch[2].l_um_iw[16] ;
 wire \top_I.branch[2].l_um_iw[170] ;
 wire \top_I.branch[2].l_um_iw[171] ;
 wire \top_I.branch[2].l_um_iw[172] ;
 wire \top_I.branch[2].l_um_iw[173] ;
 wire \top_I.branch[2].l_um_iw[174] ;
 wire \top_I.branch[2].l_um_iw[175] ;
 wire \top_I.branch[2].l_um_iw[176] ;
 wire \top_I.branch[2].l_um_iw[177] ;
 wire \top_I.branch[2].l_um_iw[178] ;
 wire \top_I.branch[2].l_um_iw[179] ;
 wire \top_I.branch[2].l_um_iw[17] ;
 wire \top_I.branch[2].l_um_iw[180] ;
 wire \top_I.branch[2].l_um_iw[181] ;
 wire \top_I.branch[2].l_um_iw[182] ;
 wire \top_I.branch[2].l_um_iw[183] ;
 wire \top_I.branch[2].l_um_iw[184] ;
 wire \top_I.branch[2].l_um_iw[185] ;
 wire \top_I.branch[2].l_um_iw[186] ;
 wire \top_I.branch[2].l_um_iw[187] ;
 wire \top_I.branch[2].l_um_iw[188] ;
 wire \top_I.branch[2].l_um_iw[189] ;
 wire \top_I.branch[2].l_um_iw[18] ;
 wire \top_I.branch[2].l_um_iw[190] ;
 wire \top_I.branch[2].l_um_iw[191] ;
 wire \top_I.branch[2].l_um_iw[192] ;
 wire \top_I.branch[2].l_um_iw[193] ;
 wire \top_I.branch[2].l_um_iw[194] ;
 wire \top_I.branch[2].l_um_iw[195] ;
 wire \top_I.branch[2].l_um_iw[196] ;
 wire \top_I.branch[2].l_um_iw[197] ;
 wire \top_I.branch[2].l_um_iw[198] ;
 wire \top_I.branch[2].l_um_iw[199] ;
 wire \top_I.branch[2].l_um_iw[19] ;
 wire \top_I.branch[2].l_um_iw[1] ;
 wire \top_I.branch[2].l_um_iw[200] ;
 wire \top_I.branch[2].l_um_iw[201] ;
 wire \top_I.branch[2].l_um_iw[202] ;
 wire \top_I.branch[2].l_um_iw[203] ;
 wire \top_I.branch[2].l_um_iw[204] ;
 wire \top_I.branch[2].l_um_iw[205] ;
 wire \top_I.branch[2].l_um_iw[206] ;
 wire \top_I.branch[2].l_um_iw[207] ;
 wire \top_I.branch[2].l_um_iw[208] ;
 wire \top_I.branch[2].l_um_iw[209] ;
 wire \top_I.branch[2].l_um_iw[20] ;
 wire \top_I.branch[2].l_um_iw[210] ;
 wire \top_I.branch[2].l_um_iw[211] ;
 wire \top_I.branch[2].l_um_iw[212] ;
 wire \top_I.branch[2].l_um_iw[213] ;
 wire \top_I.branch[2].l_um_iw[214] ;
 wire \top_I.branch[2].l_um_iw[215] ;
 wire \top_I.branch[2].l_um_iw[216] ;
 wire \top_I.branch[2].l_um_iw[217] ;
 wire \top_I.branch[2].l_um_iw[218] ;
 wire \top_I.branch[2].l_um_iw[219] ;
 wire \top_I.branch[2].l_um_iw[21] ;
 wire \top_I.branch[2].l_um_iw[220] ;
 wire \top_I.branch[2].l_um_iw[221] ;
 wire \top_I.branch[2].l_um_iw[222] ;
 wire \top_I.branch[2].l_um_iw[223] ;
 wire \top_I.branch[2].l_um_iw[224] ;
 wire \top_I.branch[2].l_um_iw[225] ;
 wire \top_I.branch[2].l_um_iw[226] ;
 wire \top_I.branch[2].l_um_iw[227] ;
 wire \top_I.branch[2].l_um_iw[228] ;
 wire \top_I.branch[2].l_um_iw[229] ;
 wire \top_I.branch[2].l_um_iw[22] ;
 wire \top_I.branch[2].l_um_iw[230] ;
 wire \top_I.branch[2].l_um_iw[231] ;
 wire \top_I.branch[2].l_um_iw[232] ;
 wire \top_I.branch[2].l_um_iw[233] ;
 wire \top_I.branch[2].l_um_iw[234] ;
 wire \top_I.branch[2].l_um_iw[235] ;
 wire \top_I.branch[2].l_um_iw[236] ;
 wire \top_I.branch[2].l_um_iw[237] ;
 wire \top_I.branch[2].l_um_iw[238] ;
 wire \top_I.branch[2].l_um_iw[239] ;
 wire \top_I.branch[2].l_um_iw[23] ;
 wire \top_I.branch[2].l_um_iw[240] ;
 wire \top_I.branch[2].l_um_iw[241] ;
 wire \top_I.branch[2].l_um_iw[242] ;
 wire \top_I.branch[2].l_um_iw[243] ;
 wire \top_I.branch[2].l_um_iw[244] ;
 wire \top_I.branch[2].l_um_iw[245] ;
 wire \top_I.branch[2].l_um_iw[246] ;
 wire \top_I.branch[2].l_um_iw[247] ;
 wire \top_I.branch[2].l_um_iw[248] ;
 wire \top_I.branch[2].l_um_iw[249] ;
 wire \top_I.branch[2].l_um_iw[24] ;
 wire \top_I.branch[2].l_um_iw[250] ;
 wire \top_I.branch[2].l_um_iw[251] ;
 wire \top_I.branch[2].l_um_iw[252] ;
 wire \top_I.branch[2].l_um_iw[253] ;
 wire \top_I.branch[2].l_um_iw[254] ;
 wire \top_I.branch[2].l_um_iw[255] ;
 wire \top_I.branch[2].l_um_iw[256] ;
 wire \top_I.branch[2].l_um_iw[257] ;
 wire \top_I.branch[2].l_um_iw[258] ;
 wire \top_I.branch[2].l_um_iw[259] ;
 wire \top_I.branch[2].l_um_iw[25] ;
 wire \top_I.branch[2].l_um_iw[260] ;
 wire \top_I.branch[2].l_um_iw[261] ;
 wire \top_I.branch[2].l_um_iw[262] ;
 wire \top_I.branch[2].l_um_iw[263] ;
 wire \top_I.branch[2].l_um_iw[264] ;
 wire \top_I.branch[2].l_um_iw[265] ;
 wire \top_I.branch[2].l_um_iw[266] ;
 wire \top_I.branch[2].l_um_iw[267] ;
 wire \top_I.branch[2].l_um_iw[268] ;
 wire \top_I.branch[2].l_um_iw[269] ;
 wire \top_I.branch[2].l_um_iw[26] ;
 wire \top_I.branch[2].l_um_iw[270] ;
 wire \top_I.branch[2].l_um_iw[271] ;
 wire \top_I.branch[2].l_um_iw[272] ;
 wire \top_I.branch[2].l_um_iw[273] ;
 wire \top_I.branch[2].l_um_iw[274] ;
 wire \top_I.branch[2].l_um_iw[275] ;
 wire \top_I.branch[2].l_um_iw[276] ;
 wire \top_I.branch[2].l_um_iw[277] ;
 wire \top_I.branch[2].l_um_iw[278] ;
 wire \top_I.branch[2].l_um_iw[279] ;
 wire \top_I.branch[2].l_um_iw[27] ;
 wire \top_I.branch[2].l_um_iw[280] ;
 wire \top_I.branch[2].l_um_iw[281] ;
 wire \top_I.branch[2].l_um_iw[282] ;
 wire \top_I.branch[2].l_um_iw[283] ;
 wire \top_I.branch[2].l_um_iw[284] ;
 wire \top_I.branch[2].l_um_iw[285] ;
 wire \top_I.branch[2].l_um_iw[286] ;
 wire \top_I.branch[2].l_um_iw[287] ;
 wire \top_I.branch[2].l_um_iw[28] ;
 wire \top_I.branch[2].l_um_iw[29] ;
 wire \top_I.branch[2].l_um_iw[2] ;
 wire \top_I.branch[2].l_um_iw[30] ;
 wire \top_I.branch[2].l_um_iw[31] ;
 wire \top_I.branch[2].l_um_iw[32] ;
 wire \top_I.branch[2].l_um_iw[33] ;
 wire \top_I.branch[2].l_um_iw[34] ;
 wire \top_I.branch[2].l_um_iw[35] ;
 wire \top_I.branch[2].l_um_iw[36] ;
 wire \top_I.branch[2].l_um_iw[37] ;
 wire \top_I.branch[2].l_um_iw[38] ;
 wire \top_I.branch[2].l_um_iw[39] ;
 wire \top_I.branch[2].l_um_iw[3] ;
 wire \top_I.branch[2].l_um_iw[40] ;
 wire \top_I.branch[2].l_um_iw[41] ;
 wire \top_I.branch[2].l_um_iw[42] ;
 wire \top_I.branch[2].l_um_iw[43] ;
 wire \top_I.branch[2].l_um_iw[44] ;
 wire \top_I.branch[2].l_um_iw[45] ;
 wire \top_I.branch[2].l_um_iw[46] ;
 wire \top_I.branch[2].l_um_iw[47] ;
 wire \top_I.branch[2].l_um_iw[48] ;
 wire \top_I.branch[2].l_um_iw[49] ;
 wire \top_I.branch[2].l_um_iw[4] ;
 wire \top_I.branch[2].l_um_iw[50] ;
 wire \top_I.branch[2].l_um_iw[51] ;
 wire \top_I.branch[2].l_um_iw[52] ;
 wire \top_I.branch[2].l_um_iw[53] ;
 wire \top_I.branch[2].l_um_iw[54] ;
 wire \top_I.branch[2].l_um_iw[55] ;
 wire \top_I.branch[2].l_um_iw[56] ;
 wire \top_I.branch[2].l_um_iw[57] ;
 wire \top_I.branch[2].l_um_iw[58] ;
 wire \top_I.branch[2].l_um_iw[59] ;
 wire \top_I.branch[2].l_um_iw[5] ;
 wire \top_I.branch[2].l_um_iw[60] ;
 wire \top_I.branch[2].l_um_iw[61] ;
 wire \top_I.branch[2].l_um_iw[62] ;
 wire \top_I.branch[2].l_um_iw[63] ;
 wire \top_I.branch[2].l_um_iw[64] ;
 wire \top_I.branch[2].l_um_iw[65] ;
 wire \top_I.branch[2].l_um_iw[66] ;
 wire \top_I.branch[2].l_um_iw[67] ;
 wire \top_I.branch[2].l_um_iw[68] ;
 wire \top_I.branch[2].l_um_iw[69] ;
 wire \top_I.branch[2].l_um_iw[6] ;
 wire \top_I.branch[2].l_um_iw[70] ;
 wire \top_I.branch[2].l_um_iw[71] ;
 wire \top_I.branch[2].l_um_iw[72] ;
 wire \top_I.branch[2].l_um_iw[73] ;
 wire \top_I.branch[2].l_um_iw[74] ;
 wire \top_I.branch[2].l_um_iw[75] ;
 wire \top_I.branch[2].l_um_iw[76] ;
 wire \top_I.branch[2].l_um_iw[77] ;
 wire \top_I.branch[2].l_um_iw[78] ;
 wire \top_I.branch[2].l_um_iw[79] ;
 wire \top_I.branch[2].l_um_iw[7] ;
 wire \top_I.branch[2].l_um_iw[80] ;
 wire \top_I.branch[2].l_um_iw[81] ;
 wire \top_I.branch[2].l_um_iw[82] ;
 wire \top_I.branch[2].l_um_iw[83] ;
 wire \top_I.branch[2].l_um_iw[84] ;
 wire \top_I.branch[2].l_um_iw[85] ;
 wire \top_I.branch[2].l_um_iw[86] ;
 wire \top_I.branch[2].l_um_iw[87] ;
 wire \top_I.branch[2].l_um_iw[88] ;
 wire \top_I.branch[2].l_um_iw[89] ;
 wire \top_I.branch[2].l_um_iw[8] ;
 wire \top_I.branch[2].l_um_iw[90] ;
 wire \top_I.branch[2].l_um_iw[91] ;
 wire \top_I.branch[2].l_um_iw[92] ;
 wire \top_I.branch[2].l_um_iw[93] ;
 wire \top_I.branch[2].l_um_iw[94] ;
 wire \top_I.branch[2].l_um_iw[95] ;
 wire \top_I.branch[2].l_um_iw[96] ;
 wire \top_I.branch[2].l_um_iw[97] ;
 wire \top_I.branch[2].l_um_iw[98] ;
 wire \top_I.branch[2].l_um_iw[99] ;
 wire \top_I.branch[2].l_um_iw[9] ;
 wire \top_I.branch[2].l_um_k_zero[0] ;
 wire \top_I.branch[2].l_um_k_zero[10] ;
 wire \top_I.branch[2].l_um_k_zero[11] ;
 wire \top_I.branch[2].l_um_k_zero[12] ;
 wire \top_I.branch[2].l_um_k_zero[13] ;
 wire \top_I.branch[2].l_um_k_zero[14] ;
 wire \top_I.branch[2].l_um_k_zero[15] ;
 wire \top_I.branch[2].l_um_k_zero[1] ;
 wire \top_I.branch[2].l_um_k_zero[2] ;
 wire \top_I.branch[2].l_um_k_zero[3] ;
 wire \top_I.branch[2].l_um_k_zero[4] ;
 wire \top_I.branch[2].l_um_k_zero[5] ;
 wire \top_I.branch[2].l_um_k_zero[6] ;
 wire \top_I.branch[2].l_um_k_zero[7] ;
 wire \top_I.branch[2].l_um_k_zero[8] ;
 wire \top_I.branch[2].l_um_k_zero[9] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[3].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[3].l_k_one ;
 wire \top_I.branch[3].l_k_zero ;
 wire \top_I.branch[3].l_um_ena[0] ;
 wire \top_I.branch[3].l_um_ena[10] ;
 wire \top_I.branch[3].l_um_ena[11] ;
 wire \top_I.branch[3].l_um_ena[12] ;
 wire \top_I.branch[3].l_um_ena[13] ;
 wire \top_I.branch[3].l_um_ena[14] ;
 wire \top_I.branch[3].l_um_ena[15] ;
 wire \top_I.branch[3].l_um_ena[1] ;
 wire \top_I.branch[3].l_um_ena[2] ;
 wire \top_I.branch[3].l_um_ena[3] ;
 wire \top_I.branch[3].l_um_ena[4] ;
 wire \top_I.branch[3].l_um_ena[5] ;
 wire \top_I.branch[3].l_um_ena[6] ;
 wire \top_I.branch[3].l_um_ena[7] ;
 wire \top_I.branch[3].l_um_ena[8] ;
 wire \top_I.branch[3].l_um_ena[9] ;
 wire \top_I.branch[3].l_um_iw[0] ;
 wire \top_I.branch[3].l_um_iw[100] ;
 wire \top_I.branch[3].l_um_iw[101] ;
 wire \top_I.branch[3].l_um_iw[102] ;
 wire \top_I.branch[3].l_um_iw[103] ;
 wire \top_I.branch[3].l_um_iw[104] ;
 wire \top_I.branch[3].l_um_iw[105] ;
 wire \top_I.branch[3].l_um_iw[106] ;
 wire \top_I.branch[3].l_um_iw[107] ;
 wire \top_I.branch[3].l_um_iw[108] ;
 wire \top_I.branch[3].l_um_iw[109] ;
 wire \top_I.branch[3].l_um_iw[10] ;
 wire \top_I.branch[3].l_um_iw[110] ;
 wire \top_I.branch[3].l_um_iw[111] ;
 wire \top_I.branch[3].l_um_iw[112] ;
 wire \top_I.branch[3].l_um_iw[113] ;
 wire \top_I.branch[3].l_um_iw[114] ;
 wire \top_I.branch[3].l_um_iw[115] ;
 wire \top_I.branch[3].l_um_iw[116] ;
 wire \top_I.branch[3].l_um_iw[117] ;
 wire \top_I.branch[3].l_um_iw[118] ;
 wire \top_I.branch[3].l_um_iw[119] ;
 wire \top_I.branch[3].l_um_iw[11] ;
 wire \top_I.branch[3].l_um_iw[120] ;
 wire \top_I.branch[3].l_um_iw[121] ;
 wire \top_I.branch[3].l_um_iw[122] ;
 wire \top_I.branch[3].l_um_iw[123] ;
 wire \top_I.branch[3].l_um_iw[124] ;
 wire \top_I.branch[3].l_um_iw[125] ;
 wire \top_I.branch[3].l_um_iw[126] ;
 wire \top_I.branch[3].l_um_iw[127] ;
 wire \top_I.branch[3].l_um_iw[128] ;
 wire \top_I.branch[3].l_um_iw[129] ;
 wire \top_I.branch[3].l_um_iw[12] ;
 wire \top_I.branch[3].l_um_iw[130] ;
 wire \top_I.branch[3].l_um_iw[131] ;
 wire \top_I.branch[3].l_um_iw[132] ;
 wire \top_I.branch[3].l_um_iw[133] ;
 wire \top_I.branch[3].l_um_iw[134] ;
 wire \top_I.branch[3].l_um_iw[135] ;
 wire \top_I.branch[3].l_um_iw[136] ;
 wire \top_I.branch[3].l_um_iw[137] ;
 wire \top_I.branch[3].l_um_iw[138] ;
 wire \top_I.branch[3].l_um_iw[139] ;
 wire \top_I.branch[3].l_um_iw[13] ;
 wire \top_I.branch[3].l_um_iw[140] ;
 wire \top_I.branch[3].l_um_iw[141] ;
 wire \top_I.branch[3].l_um_iw[142] ;
 wire \top_I.branch[3].l_um_iw[143] ;
 wire \top_I.branch[3].l_um_iw[144] ;
 wire \top_I.branch[3].l_um_iw[145] ;
 wire \top_I.branch[3].l_um_iw[146] ;
 wire \top_I.branch[3].l_um_iw[147] ;
 wire \top_I.branch[3].l_um_iw[148] ;
 wire \top_I.branch[3].l_um_iw[149] ;
 wire \top_I.branch[3].l_um_iw[14] ;
 wire \top_I.branch[3].l_um_iw[150] ;
 wire \top_I.branch[3].l_um_iw[151] ;
 wire \top_I.branch[3].l_um_iw[152] ;
 wire \top_I.branch[3].l_um_iw[153] ;
 wire \top_I.branch[3].l_um_iw[154] ;
 wire \top_I.branch[3].l_um_iw[155] ;
 wire \top_I.branch[3].l_um_iw[156] ;
 wire \top_I.branch[3].l_um_iw[157] ;
 wire \top_I.branch[3].l_um_iw[158] ;
 wire \top_I.branch[3].l_um_iw[159] ;
 wire \top_I.branch[3].l_um_iw[15] ;
 wire \top_I.branch[3].l_um_iw[160] ;
 wire \top_I.branch[3].l_um_iw[161] ;
 wire \top_I.branch[3].l_um_iw[162] ;
 wire \top_I.branch[3].l_um_iw[163] ;
 wire \top_I.branch[3].l_um_iw[164] ;
 wire \top_I.branch[3].l_um_iw[165] ;
 wire \top_I.branch[3].l_um_iw[166] ;
 wire \top_I.branch[3].l_um_iw[167] ;
 wire \top_I.branch[3].l_um_iw[168] ;
 wire \top_I.branch[3].l_um_iw[169] ;
 wire \top_I.branch[3].l_um_iw[16] ;
 wire \top_I.branch[3].l_um_iw[170] ;
 wire \top_I.branch[3].l_um_iw[171] ;
 wire \top_I.branch[3].l_um_iw[172] ;
 wire \top_I.branch[3].l_um_iw[173] ;
 wire \top_I.branch[3].l_um_iw[174] ;
 wire \top_I.branch[3].l_um_iw[175] ;
 wire \top_I.branch[3].l_um_iw[176] ;
 wire \top_I.branch[3].l_um_iw[177] ;
 wire \top_I.branch[3].l_um_iw[178] ;
 wire \top_I.branch[3].l_um_iw[179] ;
 wire \top_I.branch[3].l_um_iw[17] ;
 wire \top_I.branch[3].l_um_iw[180] ;
 wire \top_I.branch[3].l_um_iw[181] ;
 wire \top_I.branch[3].l_um_iw[182] ;
 wire \top_I.branch[3].l_um_iw[183] ;
 wire \top_I.branch[3].l_um_iw[184] ;
 wire \top_I.branch[3].l_um_iw[185] ;
 wire \top_I.branch[3].l_um_iw[186] ;
 wire \top_I.branch[3].l_um_iw[187] ;
 wire \top_I.branch[3].l_um_iw[188] ;
 wire \top_I.branch[3].l_um_iw[189] ;
 wire \top_I.branch[3].l_um_iw[18] ;
 wire \top_I.branch[3].l_um_iw[190] ;
 wire \top_I.branch[3].l_um_iw[191] ;
 wire \top_I.branch[3].l_um_iw[192] ;
 wire \top_I.branch[3].l_um_iw[193] ;
 wire \top_I.branch[3].l_um_iw[194] ;
 wire \top_I.branch[3].l_um_iw[195] ;
 wire \top_I.branch[3].l_um_iw[196] ;
 wire \top_I.branch[3].l_um_iw[197] ;
 wire \top_I.branch[3].l_um_iw[198] ;
 wire \top_I.branch[3].l_um_iw[199] ;
 wire \top_I.branch[3].l_um_iw[19] ;
 wire \top_I.branch[3].l_um_iw[1] ;
 wire \top_I.branch[3].l_um_iw[200] ;
 wire \top_I.branch[3].l_um_iw[201] ;
 wire \top_I.branch[3].l_um_iw[202] ;
 wire \top_I.branch[3].l_um_iw[203] ;
 wire \top_I.branch[3].l_um_iw[204] ;
 wire \top_I.branch[3].l_um_iw[205] ;
 wire \top_I.branch[3].l_um_iw[206] ;
 wire \top_I.branch[3].l_um_iw[207] ;
 wire \top_I.branch[3].l_um_iw[208] ;
 wire \top_I.branch[3].l_um_iw[209] ;
 wire \top_I.branch[3].l_um_iw[20] ;
 wire \top_I.branch[3].l_um_iw[210] ;
 wire \top_I.branch[3].l_um_iw[211] ;
 wire \top_I.branch[3].l_um_iw[212] ;
 wire \top_I.branch[3].l_um_iw[213] ;
 wire \top_I.branch[3].l_um_iw[214] ;
 wire \top_I.branch[3].l_um_iw[215] ;
 wire \top_I.branch[3].l_um_iw[216] ;
 wire \top_I.branch[3].l_um_iw[217] ;
 wire \top_I.branch[3].l_um_iw[218] ;
 wire \top_I.branch[3].l_um_iw[219] ;
 wire \top_I.branch[3].l_um_iw[21] ;
 wire \top_I.branch[3].l_um_iw[220] ;
 wire \top_I.branch[3].l_um_iw[221] ;
 wire \top_I.branch[3].l_um_iw[222] ;
 wire \top_I.branch[3].l_um_iw[223] ;
 wire \top_I.branch[3].l_um_iw[224] ;
 wire \top_I.branch[3].l_um_iw[225] ;
 wire \top_I.branch[3].l_um_iw[226] ;
 wire \top_I.branch[3].l_um_iw[227] ;
 wire \top_I.branch[3].l_um_iw[228] ;
 wire \top_I.branch[3].l_um_iw[229] ;
 wire \top_I.branch[3].l_um_iw[22] ;
 wire \top_I.branch[3].l_um_iw[230] ;
 wire \top_I.branch[3].l_um_iw[231] ;
 wire \top_I.branch[3].l_um_iw[232] ;
 wire \top_I.branch[3].l_um_iw[233] ;
 wire \top_I.branch[3].l_um_iw[234] ;
 wire \top_I.branch[3].l_um_iw[235] ;
 wire \top_I.branch[3].l_um_iw[236] ;
 wire \top_I.branch[3].l_um_iw[237] ;
 wire \top_I.branch[3].l_um_iw[238] ;
 wire \top_I.branch[3].l_um_iw[239] ;
 wire \top_I.branch[3].l_um_iw[23] ;
 wire \top_I.branch[3].l_um_iw[240] ;
 wire \top_I.branch[3].l_um_iw[241] ;
 wire \top_I.branch[3].l_um_iw[242] ;
 wire \top_I.branch[3].l_um_iw[243] ;
 wire \top_I.branch[3].l_um_iw[244] ;
 wire \top_I.branch[3].l_um_iw[245] ;
 wire \top_I.branch[3].l_um_iw[246] ;
 wire \top_I.branch[3].l_um_iw[247] ;
 wire \top_I.branch[3].l_um_iw[248] ;
 wire \top_I.branch[3].l_um_iw[249] ;
 wire \top_I.branch[3].l_um_iw[24] ;
 wire \top_I.branch[3].l_um_iw[250] ;
 wire \top_I.branch[3].l_um_iw[251] ;
 wire \top_I.branch[3].l_um_iw[252] ;
 wire \top_I.branch[3].l_um_iw[253] ;
 wire \top_I.branch[3].l_um_iw[254] ;
 wire \top_I.branch[3].l_um_iw[255] ;
 wire \top_I.branch[3].l_um_iw[256] ;
 wire \top_I.branch[3].l_um_iw[257] ;
 wire \top_I.branch[3].l_um_iw[258] ;
 wire \top_I.branch[3].l_um_iw[259] ;
 wire \top_I.branch[3].l_um_iw[25] ;
 wire \top_I.branch[3].l_um_iw[260] ;
 wire \top_I.branch[3].l_um_iw[261] ;
 wire \top_I.branch[3].l_um_iw[262] ;
 wire \top_I.branch[3].l_um_iw[263] ;
 wire \top_I.branch[3].l_um_iw[264] ;
 wire \top_I.branch[3].l_um_iw[265] ;
 wire \top_I.branch[3].l_um_iw[266] ;
 wire \top_I.branch[3].l_um_iw[267] ;
 wire \top_I.branch[3].l_um_iw[268] ;
 wire \top_I.branch[3].l_um_iw[269] ;
 wire \top_I.branch[3].l_um_iw[26] ;
 wire \top_I.branch[3].l_um_iw[270] ;
 wire \top_I.branch[3].l_um_iw[271] ;
 wire \top_I.branch[3].l_um_iw[272] ;
 wire \top_I.branch[3].l_um_iw[273] ;
 wire \top_I.branch[3].l_um_iw[274] ;
 wire \top_I.branch[3].l_um_iw[275] ;
 wire \top_I.branch[3].l_um_iw[276] ;
 wire \top_I.branch[3].l_um_iw[277] ;
 wire \top_I.branch[3].l_um_iw[278] ;
 wire \top_I.branch[3].l_um_iw[279] ;
 wire \top_I.branch[3].l_um_iw[27] ;
 wire \top_I.branch[3].l_um_iw[280] ;
 wire \top_I.branch[3].l_um_iw[281] ;
 wire \top_I.branch[3].l_um_iw[282] ;
 wire \top_I.branch[3].l_um_iw[283] ;
 wire \top_I.branch[3].l_um_iw[284] ;
 wire \top_I.branch[3].l_um_iw[285] ;
 wire \top_I.branch[3].l_um_iw[286] ;
 wire \top_I.branch[3].l_um_iw[287] ;
 wire \top_I.branch[3].l_um_iw[28] ;
 wire \top_I.branch[3].l_um_iw[29] ;
 wire \top_I.branch[3].l_um_iw[2] ;
 wire \top_I.branch[3].l_um_iw[30] ;
 wire \top_I.branch[3].l_um_iw[31] ;
 wire \top_I.branch[3].l_um_iw[32] ;
 wire \top_I.branch[3].l_um_iw[33] ;
 wire \top_I.branch[3].l_um_iw[34] ;
 wire \top_I.branch[3].l_um_iw[35] ;
 wire \top_I.branch[3].l_um_iw[36] ;
 wire \top_I.branch[3].l_um_iw[37] ;
 wire \top_I.branch[3].l_um_iw[38] ;
 wire \top_I.branch[3].l_um_iw[39] ;
 wire \top_I.branch[3].l_um_iw[3] ;
 wire \top_I.branch[3].l_um_iw[40] ;
 wire \top_I.branch[3].l_um_iw[41] ;
 wire \top_I.branch[3].l_um_iw[42] ;
 wire \top_I.branch[3].l_um_iw[43] ;
 wire \top_I.branch[3].l_um_iw[44] ;
 wire \top_I.branch[3].l_um_iw[45] ;
 wire \top_I.branch[3].l_um_iw[46] ;
 wire \top_I.branch[3].l_um_iw[47] ;
 wire \top_I.branch[3].l_um_iw[48] ;
 wire \top_I.branch[3].l_um_iw[49] ;
 wire \top_I.branch[3].l_um_iw[4] ;
 wire \top_I.branch[3].l_um_iw[50] ;
 wire \top_I.branch[3].l_um_iw[51] ;
 wire \top_I.branch[3].l_um_iw[52] ;
 wire \top_I.branch[3].l_um_iw[53] ;
 wire \top_I.branch[3].l_um_iw[54] ;
 wire \top_I.branch[3].l_um_iw[55] ;
 wire \top_I.branch[3].l_um_iw[56] ;
 wire \top_I.branch[3].l_um_iw[57] ;
 wire \top_I.branch[3].l_um_iw[58] ;
 wire \top_I.branch[3].l_um_iw[59] ;
 wire \top_I.branch[3].l_um_iw[5] ;
 wire \top_I.branch[3].l_um_iw[60] ;
 wire \top_I.branch[3].l_um_iw[61] ;
 wire \top_I.branch[3].l_um_iw[62] ;
 wire \top_I.branch[3].l_um_iw[63] ;
 wire \top_I.branch[3].l_um_iw[64] ;
 wire \top_I.branch[3].l_um_iw[65] ;
 wire \top_I.branch[3].l_um_iw[66] ;
 wire \top_I.branch[3].l_um_iw[67] ;
 wire \top_I.branch[3].l_um_iw[68] ;
 wire \top_I.branch[3].l_um_iw[69] ;
 wire \top_I.branch[3].l_um_iw[6] ;
 wire \top_I.branch[3].l_um_iw[70] ;
 wire \top_I.branch[3].l_um_iw[71] ;
 wire \top_I.branch[3].l_um_iw[72] ;
 wire \top_I.branch[3].l_um_iw[73] ;
 wire \top_I.branch[3].l_um_iw[74] ;
 wire \top_I.branch[3].l_um_iw[75] ;
 wire \top_I.branch[3].l_um_iw[76] ;
 wire \top_I.branch[3].l_um_iw[77] ;
 wire \top_I.branch[3].l_um_iw[78] ;
 wire \top_I.branch[3].l_um_iw[79] ;
 wire \top_I.branch[3].l_um_iw[7] ;
 wire \top_I.branch[3].l_um_iw[80] ;
 wire \top_I.branch[3].l_um_iw[81] ;
 wire \top_I.branch[3].l_um_iw[82] ;
 wire \top_I.branch[3].l_um_iw[83] ;
 wire \top_I.branch[3].l_um_iw[84] ;
 wire \top_I.branch[3].l_um_iw[85] ;
 wire \top_I.branch[3].l_um_iw[86] ;
 wire \top_I.branch[3].l_um_iw[87] ;
 wire \top_I.branch[3].l_um_iw[88] ;
 wire \top_I.branch[3].l_um_iw[89] ;
 wire \top_I.branch[3].l_um_iw[8] ;
 wire \top_I.branch[3].l_um_iw[90] ;
 wire \top_I.branch[3].l_um_iw[91] ;
 wire \top_I.branch[3].l_um_iw[92] ;
 wire \top_I.branch[3].l_um_iw[93] ;
 wire \top_I.branch[3].l_um_iw[94] ;
 wire \top_I.branch[3].l_um_iw[95] ;
 wire \top_I.branch[3].l_um_iw[96] ;
 wire \top_I.branch[3].l_um_iw[97] ;
 wire \top_I.branch[3].l_um_iw[98] ;
 wire \top_I.branch[3].l_um_iw[99] ;
 wire \top_I.branch[3].l_um_iw[9] ;
 wire \top_I.branch[3].l_um_k_zero[0] ;
 wire \top_I.branch[3].l_um_k_zero[10] ;
 wire \top_I.branch[3].l_um_k_zero[11] ;
 wire \top_I.branch[3].l_um_k_zero[12] ;
 wire \top_I.branch[3].l_um_k_zero[13] ;
 wire \top_I.branch[3].l_um_k_zero[14] ;
 wire \top_I.branch[3].l_um_k_zero[15] ;
 wire \top_I.branch[3].l_um_k_zero[1] ;
 wire \top_I.branch[3].l_um_k_zero[2] ;
 wire \top_I.branch[3].l_um_k_zero[3] ;
 wire \top_I.branch[3].l_um_k_zero[4] ;
 wire \top_I.branch[3].l_um_k_zero[5] ;
 wire \top_I.branch[3].l_um_k_zero[6] ;
 wire \top_I.branch[3].l_um_k_zero[7] ;
 wire \top_I.branch[3].l_um_k_zero[8] ;
 wire \top_I.branch[3].l_um_k_zero[9] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[4].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[0] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[1] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[2] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[3] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[4] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[5] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[6] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_oe[7] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[0] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[1] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[2] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[3] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[4] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[5] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[6] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uio_out[7] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[0] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[1] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[2] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[3] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[4] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[5] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[6] ;
 wire \top_I.branch[4].col_um[2].um_top_I.uo_out[7] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[0] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[1] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[2] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[3] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[4] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[5] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[6] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_oe[7] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[0] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[1] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[2] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[3] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[4] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[5] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[6] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uio_out[7] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[0] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[1] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[2] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[3] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[4] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[5] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[6] ;
 wire \top_I.branch[4].col_um[4].um_top_I.uo_out[7] ;
 wire \top_I.branch[4].l_k_one ;
 wire \top_I.branch[4].l_k_zero ;
 wire \top_I.branch[4].l_um_ena[0] ;
 wire \top_I.branch[4].l_um_ena[10] ;
 wire \top_I.branch[4].l_um_ena[11] ;
 wire \top_I.branch[4].l_um_ena[12] ;
 wire \top_I.branch[4].l_um_ena[13] ;
 wire \top_I.branch[4].l_um_ena[14] ;
 wire \top_I.branch[4].l_um_ena[15] ;
 wire \top_I.branch[4].l_um_ena[1] ;
 wire \top_I.branch[4].l_um_ena[2] ;
 wire \top_I.branch[4].l_um_ena[3] ;
 wire \top_I.branch[4].l_um_ena[4] ;
 wire \top_I.branch[4].l_um_ena[5] ;
 wire \top_I.branch[4].l_um_ena[6] ;
 wire \top_I.branch[4].l_um_ena[7] ;
 wire \top_I.branch[4].l_um_ena[8] ;
 wire \top_I.branch[4].l_um_ena[9] ;
 wire \top_I.branch[4].l_um_iw[0] ;
 wire \top_I.branch[4].l_um_iw[100] ;
 wire \top_I.branch[4].l_um_iw[101] ;
 wire \top_I.branch[4].l_um_iw[102] ;
 wire \top_I.branch[4].l_um_iw[103] ;
 wire \top_I.branch[4].l_um_iw[104] ;
 wire \top_I.branch[4].l_um_iw[105] ;
 wire \top_I.branch[4].l_um_iw[106] ;
 wire \top_I.branch[4].l_um_iw[107] ;
 wire \top_I.branch[4].l_um_iw[108] ;
 wire \top_I.branch[4].l_um_iw[109] ;
 wire \top_I.branch[4].l_um_iw[10] ;
 wire \top_I.branch[4].l_um_iw[110] ;
 wire \top_I.branch[4].l_um_iw[111] ;
 wire \top_I.branch[4].l_um_iw[112] ;
 wire \top_I.branch[4].l_um_iw[113] ;
 wire \top_I.branch[4].l_um_iw[114] ;
 wire \top_I.branch[4].l_um_iw[115] ;
 wire \top_I.branch[4].l_um_iw[116] ;
 wire \top_I.branch[4].l_um_iw[117] ;
 wire \top_I.branch[4].l_um_iw[118] ;
 wire \top_I.branch[4].l_um_iw[119] ;
 wire \top_I.branch[4].l_um_iw[11] ;
 wire \top_I.branch[4].l_um_iw[120] ;
 wire \top_I.branch[4].l_um_iw[121] ;
 wire \top_I.branch[4].l_um_iw[122] ;
 wire \top_I.branch[4].l_um_iw[123] ;
 wire \top_I.branch[4].l_um_iw[124] ;
 wire \top_I.branch[4].l_um_iw[125] ;
 wire \top_I.branch[4].l_um_iw[126] ;
 wire \top_I.branch[4].l_um_iw[127] ;
 wire \top_I.branch[4].l_um_iw[128] ;
 wire \top_I.branch[4].l_um_iw[129] ;
 wire \top_I.branch[4].l_um_iw[12] ;
 wire \top_I.branch[4].l_um_iw[130] ;
 wire \top_I.branch[4].l_um_iw[131] ;
 wire \top_I.branch[4].l_um_iw[132] ;
 wire \top_I.branch[4].l_um_iw[133] ;
 wire \top_I.branch[4].l_um_iw[134] ;
 wire \top_I.branch[4].l_um_iw[135] ;
 wire \top_I.branch[4].l_um_iw[136] ;
 wire \top_I.branch[4].l_um_iw[137] ;
 wire \top_I.branch[4].l_um_iw[138] ;
 wire \top_I.branch[4].l_um_iw[139] ;
 wire \top_I.branch[4].l_um_iw[13] ;
 wire \top_I.branch[4].l_um_iw[140] ;
 wire \top_I.branch[4].l_um_iw[141] ;
 wire \top_I.branch[4].l_um_iw[142] ;
 wire \top_I.branch[4].l_um_iw[143] ;
 wire \top_I.branch[4].l_um_iw[144] ;
 wire \top_I.branch[4].l_um_iw[145] ;
 wire \top_I.branch[4].l_um_iw[146] ;
 wire \top_I.branch[4].l_um_iw[147] ;
 wire \top_I.branch[4].l_um_iw[148] ;
 wire \top_I.branch[4].l_um_iw[149] ;
 wire \top_I.branch[4].l_um_iw[14] ;
 wire \top_I.branch[4].l_um_iw[150] ;
 wire \top_I.branch[4].l_um_iw[151] ;
 wire \top_I.branch[4].l_um_iw[152] ;
 wire \top_I.branch[4].l_um_iw[153] ;
 wire \top_I.branch[4].l_um_iw[154] ;
 wire \top_I.branch[4].l_um_iw[155] ;
 wire \top_I.branch[4].l_um_iw[156] ;
 wire \top_I.branch[4].l_um_iw[157] ;
 wire \top_I.branch[4].l_um_iw[158] ;
 wire \top_I.branch[4].l_um_iw[159] ;
 wire \top_I.branch[4].l_um_iw[15] ;
 wire \top_I.branch[4].l_um_iw[160] ;
 wire \top_I.branch[4].l_um_iw[161] ;
 wire \top_I.branch[4].l_um_iw[162] ;
 wire \top_I.branch[4].l_um_iw[163] ;
 wire \top_I.branch[4].l_um_iw[164] ;
 wire \top_I.branch[4].l_um_iw[165] ;
 wire \top_I.branch[4].l_um_iw[166] ;
 wire \top_I.branch[4].l_um_iw[167] ;
 wire \top_I.branch[4].l_um_iw[168] ;
 wire \top_I.branch[4].l_um_iw[169] ;
 wire \top_I.branch[4].l_um_iw[16] ;
 wire \top_I.branch[4].l_um_iw[170] ;
 wire \top_I.branch[4].l_um_iw[171] ;
 wire \top_I.branch[4].l_um_iw[172] ;
 wire \top_I.branch[4].l_um_iw[173] ;
 wire \top_I.branch[4].l_um_iw[174] ;
 wire \top_I.branch[4].l_um_iw[175] ;
 wire \top_I.branch[4].l_um_iw[176] ;
 wire \top_I.branch[4].l_um_iw[177] ;
 wire \top_I.branch[4].l_um_iw[178] ;
 wire \top_I.branch[4].l_um_iw[179] ;
 wire \top_I.branch[4].l_um_iw[17] ;
 wire \top_I.branch[4].l_um_iw[180] ;
 wire \top_I.branch[4].l_um_iw[181] ;
 wire \top_I.branch[4].l_um_iw[182] ;
 wire \top_I.branch[4].l_um_iw[183] ;
 wire \top_I.branch[4].l_um_iw[184] ;
 wire \top_I.branch[4].l_um_iw[185] ;
 wire \top_I.branch[4].l_um_iw[186] ;
 wire \top_I.branch[4].l_um_iw[187] ;
 wire \top_I.branch[4].l_um_iw[188] ;
 wire \top_I.branch[4].l_um_iw[189] ;
 wire \top_I.branch[4].l_um_iw[18] ;
 wire \top_I.branch[4].l_um_iw[190] ;
 wire \top_I.branch[4].l_um_iw[191] ;
 wire \top_I.branch[4].l_um_iw[192] ;
 wire \top_I.branch[4].l_um_iw[193] ;
 wire \top_I.branch[4].l_um_iw[194] ;
 wire \top_I.branch[4].l_um_iw[195] ;
 wire \top_I.branch[4].l_um_iw[196] ;
 wire \top_I.branch[4].l_um_iw[197] ;
 wire \top_I.branch[4].l_um_iw[198] ;
 wire \top_I.branch[4].l_um_iw[199] ;
 wire \top_I.branch[4].l_um_iw[19] ;
 wire \top_I.branch[4].l_um_iw[1] ;
 wire \top_I.branch[4].l_um_iw[200] ;
 wire \top_I.branch[4].l_um_iw[201] ;
 wire \top_I.branch[4].l_um_iw[202] ;
 wire \top_I.branch[4].l_um_iw[203] ;
 wire \top_I.branch[4].l_um_iw[204] ;
 wire \top_I.branch[4].l_um_iw[205] ;
 wire \top_I.branch[4].l_um_iw[206] ;
 wire \top_I.branch[4].l_um_iw[207] ;
 wire \top_I.branch[4].l_um_iw[208] ;
 wire \top_I.branch[4].l_um_iw[209] ;
 wire \top_I.branch[4].l_um_iw[20] ;
 wire \top_I.branch[4].l_um_iw[210] ;
 wire \top_I.branch[4].l_um_iw[211] ;
 wire \top_I.branch[4].l_um_iw[212] ;
 wire \top_I.branch[4].l_um_iw[213] ;
 wire \top_I.branch[4].l_um_iw[214] ;
 wire \top_I.branch[4].l_um_iw[215] ;
 wire \top_I.branch[4].l_um_iw[216] ;
 wire \top_I.branch[4].l_um_iw[217] ;
 wire \top_I.branch[4].l_um_iw[218] ;
 wire \top_I.branch[4].l_um_iw[219] ;
 wire \top_I.branch[4].l_um_iw[21] ;
 wire \top_I.branch[4].l_um_iw[220] ;
 wire \top_I.branch[4].l_um_iw[221] ;
 wire \top_I.branch[4].l_um_iw[222] ;
 wire \top_I.branch[4].l_um_iw[223] ;
 wire \top_I.branch[4].l_um_iw[224] ;
 wire \top_I.branch[4].l_um_iw[225] ;
 wire \top_I.branch[4].l_um_iw[226] ;
 wire \top_I.branch[4].l_um_iw[227] ;
 wire \top_I.branch[4].l_um_iw[228] ;
 wire \top_I.branch[4].l_um_iw[229] ;
 wire \top_I.branch[4].l_um_iw[22] ;
 wire \top_I.branch[4].l_um_iw[230] ;
 wire \top_I.branch[4].l_um_iw[231] ;
 wire \top_I.branch[4].l_um_iw[232] ;
 wire \top_I.branch[4].l_um_iw[233] ;
 wire \top_I.branch[4].l_um_iw[234] ;
 wire \top_I.branch[4].l_um_iw[235] ;
 wire \top_I.branch[4].l_um_iw[236] ;
 wire \top_I.branch[4].l_um_iw[237] ;
 wire \top_I.branch[4].l_um_iw[238] ;
 wire \top_I.branch[4].l_um_iw[239] ;
 wire \top_I.branch[4].l_um_iw[23] ;
 wire \top_I.branch[4].l_um_iw[240] ;
 wire \top_I.branch[4].l_um_iw[241] ;
 wire \top_I.branch[4].l_um_iw[242] ;
 wire \top_I.branch[4].l_um_iw[243] ;
 wire \top_I.branch[4].l_um_iw[244] ;
 wire \top_I.branch[4].l_um_iw[245] ;
 wire \top_I.branch[4].l_um_iw[246] ;
 wire \top_I.branch[4].l_um_iw[247] ;
 wire \top_I.branch[4].l_um_iw[248] ;
 wire \top_I.branch[4].l_um_iw[249] ;
 wire \top_I.branch[4].l_um_iw[24] ;
 wire \top_I.branch[4].l_um_iw[250] ;
 wire \top_I.branch[4].l_um_iw[251] ;
 wire \top_I.branch[4].l_um_iw[252] ;
 wire \top_I.branch[4].l_um_iw[253] ;
 wire \top_I.branch[4].l_um_iw[254] ;
 wire \top_I.branch[4].l_um_iw[255] ;
 wire \top_I.branch[4].l_um_iw[256] ;
 wire \top_I.branch[4].l_um_iw[257] ;
 wire \top_I.branch[4].l_um_iw[258] ;
 wire \top_I.branch[4].l_um_iw[259] ;
 wire \top_I.branch[4].l_um_iw[25] ;
 wire \top_I.branch[4].l_um_iw[260] ;
 wire \top_I.branch[4].l_um_iw[261] ;
 wire \top_I.branch[4].l_um_iw[262] ;
 wire \top_I.branch[4].l_um_iw[263] ;
 wire \top_I.branch[4].l_um_iw[264] ;
 wire \top_I.branch[4].l_um_iw[265] ;
 wire \top_I.branch[4].l_um_iw[266] ;
 wire \top_I.branch[4].l_um_iw[267] ;
 wire \top_I.branch[4].l_um_iw[268] ;
 wire \top_I.branch[4].l_um_iw[269] ;
 wire \top_I.branch[4].l_um_iw[26] ;
 wire \top_I.branch[4].l_um_iw[270] ;
 wire \top_I.branch[4].l_um_iw[271] ;
 wire \top_I.branch[4].l_um_iw[272] ;
 wire \top_I.branch[4].l_um_iw[273] ;
 wire \top_I.branch[4].l_um_iw[274] ;
 wire \top_I.branch[4].l_um_iw[275] ;
 wire \top_I.branch[4].l_um_iw[276] ;
 wire \top_I.branch[4].l_um_iw[277] ;
 wire \top_I.branch[4].l_um_iw[278] ;
 wire \top_I.branch[4].l_um_iw[279] ;
 wire \top_I.branch[4].l_um_iw[27] ;
 wire \top_I.branch[4].l_um_iw[280] ;
 wire \top_I.branch[4].l_um_iw[281] ;
 wire \top_I.branch[4].l_um_iw[282] ;
 wire \top_I.branch[4].l_um_iw[283] ;
 wire \top_I.branch[4].l_um_iw[284] ;
 wire \top_I.branch[4].l_um_iw[285] ;
 wire \top_I.branch[4].l_um_iw[286] ;
 wire \top_I.branch[4].l_um_iw[287] ;
 wire \top_I.branch[4].l_um_iw[28] ;
 wire \top_I.branch[4].l_um_iw[29] ;
 wire \top_I.branch[4].l_um_iw[2] ;
 wire \top_I.branch[4].l_um_iw[30] ;
 wire \top_I.branch[4].l_um_iw[31] ;
 wire \top_I.branch[4].l_um_iw[32] ;
 wire \top_I.branch[4].l_um_iw[33] ;
 wire \top_I.branch[4].l_um_iw[34] ;
 wire \top_I.branch[4].l_um_iw[35] ;
 wire \top_I.branch[4].l_um_iw[36] ;
 wire \top_I.branch[4].l_um_iw[37] ;
 wire \top_I.branch[4].l_um_iw[38] ;
 wire \top_I.branch[4].l_um_iw[39] ;
 wire \top_I.branch[4].l_um_iw[3] ;
 wire \top_I.branch[4].l_um_iw[40] ;
 wire \top_I.branch[4].l_um_iw[41] ;
 wire \top_I.branch[4].l_um_iw[42] ;
 wire \top_I.branch[4].l_um_iw[43] ;
 wire \top_I.branch[4].l_um_iw[44] ;
 wire \top_I.branch[4].l_um_iw[45] ;
 wire \top_I.branch[4].l_um_iw[46] ;
 wire \top_I.branch[4].l_um_iw[47] ;
 wire \top_I.branch[4].l_um_iw[48] ;
 wire \top_I.branch[4].l_um_iw[49] ;
 wire \top_I.branch[4].l_um_iw[4] ;
 wire \top_I.branch[4].l_um_iw[50] ;
 wire \top_I.branch[4].l_um_iw[51] ;
 wire \top_I.branch[4].l_um_iw[52] ;
 wire \top_I.branch[4].l_um_iw[53] ;
 wire \top_I.branch[4].l_um_iw[54] ;
 wire \top_I.branch[4].l_um_iw[55] ;
 wire \top_I.branch[4].l_um_iw[56] ;
 wire \top_I.branch[4].l_um_iw[57] ;
 wire \top_I.branch[4].l_um_iw[58] ;
 wire \top_I.branch[4].l_um_iw[59] ;
 wire \top_I.branch[4].l_um_iw[5] ;
 wire \top_I.branch[4].l_um_iw[60] ;
 wire \top_I.branch[4].l_um_iw[61] ;
 wire \top_I.branch[4].l_um_iw[62] ;
 wire \top_I.branch[4].l_um_iw[63] ;
 wire \top_I.branch[4].l_um_iw[64] ;
 wire \top_I.branch[4].l_um_iw[65] ;
 wire \top_I.branch[4].l_um_iw[66] ;
 wire \top_I.branch[4].l_um_iw[67] ;
 wire \top_I.branch[4].l_um_iw[68] ;
 wire \top_I.branch[4].l_um_iw[69] ;
 wire \top_I.branch[4].l_um_iw[6] ;
 wire \top_I.branch[4].l_um_iw[70] ;
 wire \top_I.branch[4].l_um_iw[71] ;
 wire \top_I.branch[4].l_um_iw[72] ;
 wire \top_I.branch[4].l_um_iw[73] ;
 wire \top_I.branch[4].l_um_iw[74] ;
 wire \top_I.branch[4].l_um_iw[75] ;
 wire \top_I.branch[4].l_um_iw[76] ;
 wire \top_I.branch[4].l_um_iw[77] ;
 wire \top_I.branch[4].l_um_iw[78] ;
 wire \top_I.branch[4].l_um_iw[79] ;
 wire \top_I.branch[4].l_um_iw[7] ;
 wire \top_I.branch[4].l_um_iw[80] ;
 wire \top_I.branch[4].l_um_iw[81] ;
 wire \top_I.branch[4].l_um_iw[82] ;
 wire \top_I.branch[4].l_um_iw[83] ;
 wire \top_I.branch[4].l_um_iw[84] ;
 wire \top_I.branch[4].l_um_iw[85] ;
 wire \top_I.branch[4].l_um_iw[86] ;
 wire \top_I.branch[4].l_um_iw[87] ;
 wire \top_I.branch[4].l_um_iw[88] ;
 wire \top_I.branch[4].l_um_iw[89] ;
 wire \top_I.branch[4].l_um_iw[8] ;
 wire \top_I.branch[4].l_um_iw[90] ;
 wire \top_I.branch[4].l_um_iw[91] ;
 wire \top_I.branch[4].l_um_iw[92] ;
 wire \top_I.branch[4].l_um_iw[93] ;
 wire \top_I.branch[4].l_um_iw[94] ;
 wire \top_I.branch[4].l_um_iw[95] ;
 wire \top_I.branch[4].l_um_iw[96] ;
 wire \top_I.branch[4].l_um_iw[97] ;
 wire \top_I.branch[4].l_um_iw[98] ;
 wire \top_I.branch[4].l_um_iw[99] ;
 wire \top_I.branch[4].l_um_iw[9] ;
 wire \top_I.branch[4].l_um_k_zero[0] ;
 wire \top_I.branch[4].l_um_k_zero[10] ;
 wire \top_I.branch[4].l_um_k_zero[11] ;
 wire \top_I.branch[4].l_um_k_zero[12] ;
 wire \top_I.branch[4].l_um_k_zero[13] ;
 wire \top_I.branch[4].l_um_k_zero[14] ;
 wire \top_I.branch[4].l_um_k_zero[15] ;
 wire \top_I.branch[4].l_um_k_zero[1] ;
 wire \top_I.branch[4].l_um_k_zero[2] ;
 wire \top_I.branch[4].l_um_k_zero[3] ;
 wire \top_I.branch[4].l_um_k_zero[4] ;
 wire \top_I.branch[4].l_um_k_zero[5] ;
 wire \top_I.branch[4].l_um_k_zero[6] ;
 wire \top_I.branch[4].l_um_k_zero[7] ;
 wire \top_I.branch[4].l_um_k_zero[8] ;
 wire \top_I.branch[4].l_um_k_zero[9] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[5].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[5].l_k_one ;
 wire \top_I.branch[5].l_k_zero ;
 wire \top_I.branch[5].l_um_ena[0] ;
 wire \top_I.branch[5].l_um_ena[10] ;
 wire \top_I.branch[5].l_um_ena[11] ;
 wire \top_I.branch[5].l_um_ena[12] ;
 wire \top_I.branch[5].l_um_ena[13] ;
 wire \top_I.branch[5].l_um_ena[14] ;
 wire \top_I.branch[5].l_um_ena[15] ;
 wire \top_I.branch[5].l_um_ena[1] ;
 wire \top_I.branch[5].l_um_ena[2] ;
 wire \top_I.branch[5].l_um_ena[3] ;
 wire \top_I.branch[5].l_um_ena[4] ;
 wire \top_I.branch[5].l_um_ena[5] ;
 wire \top_I.branch[5].l_um_ena[6] ;
 wire \top_I.branch[5].l_um_ena[7] ;
 wire \top_I.branch[5].l_um_ena[8] ;
 wire \top_I.branch[5].l_um_ena[9] ;
 wire \top_I.branch[5].l_um_iw[0] ;
 wire \top_I.branch[5].l_um_iw[100] ;
 wire \top_I.branch[5].l_um_iw[101] ;
 wire \top_I.branch[5].l_um_iw[102] ;
 wire \top_I.branch[5].l_um_iw[103] ;
 wire \top_I.branch[5].l_um_iw[104] ;
 wire \top_I.branch[5].l_um_iw[105] ;
 wire \top_I.branch[5].l_um_iw[106] ;
 wire \top_I.branch[5].l_um_iw[107] ;
 wire \top_I.branch[5].l_um_iw[108] ;
 wire \top_I.branch[5].l_um_iw[109] ;
 wire \top_I.branch[5].l_um_iw[10] ;
 wire \top_I.branch[5].l_um_iw[110] ;
 wire \top_I.branch[5].l_um_iw[111] ;
 wire \top_I.branch[5].l_um_iw[112] ;
 wire \top_I.branch[5].l_um_iw[113] ;
 wire \top_I.branch[5].l_um_iw[114] ;
 wire \top_I.branch[5].l_um_iw[115] ;
 wire \top_I.branch[5].l_um_iw[116] ;
 wire \top_I.branch[5].l_um_iw[117] ;
 wire \top_I.branch[5].l_um_iw[118] ;
 wire \top_I.branch[5].l_um_iw[119] ;
 wire \top_I.branch[5].l_um_iw[11] ;
 wire \top_I.branch[5].l_um_iw[120] ;
 wire \top_I.branch[5].l_um_iw[121] ;
 wire \top_I.branch[5].l_um_iw[122] ;
 wire \top_I.branch[5].l_um_iw[123] ;
 wire \top_I.branch[5].l_um_iw[124] ;
 wire \top_I.branch[5].l_um_iw[125] ;
 wire \top_I.branch[5].l_um_iw[126] ;
 wire \top_I.branch[5].l_um_iw[127] ;
 wire \top_I.branch[5].l_um_iw[128] ;
 wire \top_I.branch[5].l_um_iw[129] ;
 wire \top_I.branch[5].l_um_iw[12] ;
 wire \top_I.branch[5].l_um_iw[130] ;
 wire \top_I.branch[5].l_um_iw[131] ;
 wire \top_I.branch[5].l_um_iw[132] ;
 wire \top_I.branch[5].l_um_iw[133] ;
 wire \top_I.branch[5].l_um_iw[134] ;
 wire \top_I.branch[5].l_um_iw[135] ;
 wire \top_I.branch[5].l_um_iw[136] ;
 wire \top_I.branch[5].l_um_iw[137] ;
 wire \top_I.branch[5].l_um_iw[138] ;
 wire \top_I.branch[5].l_um_iw[139] ;
 wire \top_I.branch[5].l_um_iw[13] ;
 wire \top_I.branch[5].l_um_iw[140] ;
 wire \top_I.branch[5].l_um_iw[141] ;
 wire \top_I.branch[5].l_um_iw[142] ;
 wire \top_I.branch[5].l_um_iw[143] ;
 wire \top_I.branch[5].l_um_iw[144] ;
 wire \top_I.branch[5].l_um_iw[145] ;
 wire \top_I.branch[5].l_um_iw[146] ;
 wire \top_I.branch[5].l_um_iw[147] ;
 wire \top_I.branch[5].l_um_iw[148] ;
 wire \top_I.branch[5].l_um_iw[149] ;
 wire \top_I.branch[5].l_um_iw[14] ;
 wire \top_I.branch[5].l_um_iw[150] ;
 wire \top_I.branch[5].l_um_iw[151] ;
 wire \top_I.branch[5].l_um_iw[152] ;
 wire \top_I.branch[5].l_um_iw[153] ;
 wire \top_I.branch[5].l_um_iw[154] ;
 wire \top_I.branch[5].l_um_iw[155] ;
 wire \top_I.branch[5].l_um_iw[156] ;
 wire \top_I.branch[5].l_um_iw[157] ;
 wire \top_I.branch[5].l_um_iw[158] ;
 wire \top_I.branch[5].l_um_iw[159] ;
 wire \top_I.branch[5].l_um_iw[15] ;
 wire \top_I.branch[5].l_um_iw[160] ;
 wire \top_I.branch[5].l_um_iw[161] ;
 wire \top_I.branch[5].l_um_iw[162] ;
 wire \top_I.branch[5].l_um_iw[163] ;
 wire \top_I.branch[5].l_um_iw[164] ;
 wire \top_I.branch[5].l_um_iw[165] ;
 wire \top_I.branch[5].l_um_iw[166] ;
 wire \top_I.branch[5].l_um_iw[167] ;
 wire \top_I.branch[5].l_um_iw[168] ;
 wire \top_I.branch[5].l_um_iw[169] ;
 wire \top_I.branch[5].l_um_iw[16] ;
 wire \top_I.branch[5].l_um_iw[170] ;
 wire \top_I.branch[5].l_um_iw[171] ;
 wire \top_I.branch[5].l_um_iw[172] ;
 wire \top_I.branch[5].l_um_iw[173] ;
 wire \top_I.branch[5].l_um_iw[174] ;
 wire \top_I.branch[5].l_um_iw[175] ;
 wire \top_I.branch[5].l_um_iw[176] ;
 wire \top_I.branch[5].l_um_iw[177] ;
 wire \top_I.branch[5].l_um_iw[178] ;
 wire \top_I.branch[5].l_um_iw[179] ;
 wire \top_I.branch[5].l_um_iw[17] ;
 wire \top_I.branch[5].l_um_iw[180] ;
 wire \top_I.branch[5].l_um_iw[181] ;
 wire \top_I.branch[5].l_um_iw[182] ;
 wire \top_I.branch[5].l_um_iw[183] ;
 wire \top_I.branch[5].l_um_iw[184] ;
 wire \top_I.branch[5].l_um_iw[185] ;
 wire \top_I.branch[5].l_um_iw[186] ;
 wire \top_I.branch[5].l_um_iw[187] ;
 wire \top_I.branch[5].l_um_iw[188] ;
 wire \top_I.branch[5].l_um_iw[189] ;
 wire \top_I.branch[5].l_um_iw[18] ;
 wire \top_I.branch[5].l_um_iw[190] ;
 wire \top_I.branch[5].l_um_iw[191] ;
 wire \top_I.branch[5].l_um_iw[192] ;
 wire \top_I.branch[5].l_um_iw[193] ;
 wire \top_I.branch[5].l_um_iw[194] ;
 wire \top_I.branch[5].l_um_iw[195] ;
 wire \top_I.branch[5].l_um_iw[196] ;
 wire \top_I.branch[5].l_um_iw[197] ;
 wire \top_I.branch[5].l_um_iw[198] ;
 wire \top_I.branch[5].l_um_iw[199] ;
 wire \top_I.branch[5].l_um_iw[19] ;
 wire \top_I.branch[5].l_um_iw[1] ;
 wire \top_I.branch[5].l_um_iw[200] ;
 wire \top_I.branch[5].l_um_iw[201] ;
 wire \top_I.branch[5].l_um_iw[202] ;
 wire \top_I.branch[5].l_um_iw[203] ;
 wire \top_I.branch[5].l_um_iw[204] ;
 wire \top_I.branch[5].l_um_iw[205] ;
 wire \top_I.branch[5].l_um_iw[206] ;
 wire \top_I.branch[5].l_um_iw[207] ;
 wire \top_I.branch[5].l_um_iw[208] ;
 wire \top_I.branch[5].l_um_iw[209] ;
 wire \top_I.branch[5].l_um_iw[20] ;
 wire \top_I.branch[5].l_um_iw[210] ;
 wire \top_I.branch[5].l_um_iw[211] ;
 wire \top_I.branch[5].l_um_iw[212] ;
 wire \top_I.branch[5].l_um_iw[213] ;
 wire \top_I.branch[5].l_um_iw[214] ;
 wire \top_I.branch[5].l_um_iw[215] ;
 wire \top_I.branch[5].l_um_iw[216] ;
 wire \top_I.branch[5].l_um_iw[217] ;
 wire \top_I.branch[5].l_um_iw[218] ;
 wire \top_I.branch[5].l_um_iw[219] ;
 wire \top_I.branch[5].l_um_iw[21] ;
 wire \top_I.branch[5].l_um_iw[220] ;
 wire \top_I.branch[5].l_um_iw[221] ;
 wire \top_I.branch[5].l_um_iw[222] ;
 wire \top_I.branch[5].l_um_iw[223] ;
 wire \top_I.branch[5].l_um_iw[224] ;
 wire \top_I.branch[5].l_um_iw[225] ;
 wire \top_I.branch[5].l_um_iw[226] ;
 wire \top_I.branch[5].l_um_iw[227] ;
 wire \top_I.branch[5].l_um_iw[228] ;
 wire \top_I.branch[5].l_um_iw[229] ;
 wire \top_I.branch[5].l_um_iw[22] ;
 wire \top_I.branch[5].l_um_iw[230] ;
 wire \top_I.branch[5].l_um_iw[231] ;
 wire \top_I.branch[5].l_um_iw[232] ;
 wire \top_I.branch[5].l_um_iw[233] ;
 wire \top_I.branch[5].l_um_iw[234] ;
 wire \top_I.branch[5].l_um_iw[235] ;
 wire \top_I.branch[5].l_um_iw[236] ;
 wire \top_I.branch[5].l_um_iw[237] ;
 wire \top_I.branch[5].l_um_iw[238] ;
 wire \top_I.branch[5].l_um_iw[239] ;
 wire \top_I.branch[5].l_um_iw[23] ;
 wire \top_I.branch[5].l_um_iw[240] ;
 wire \top_I.branch[5].l_um_iw[241] ;
 wire \top_I.branch[5].l_um_iw[242] ;
 wire \top_I.branch[5].l_um_iw[243] ;
 wire \top_I.branch[5].l_um_iw[244] ;
 wire \top_I.branch[5].l_um_iw[245] ;
 wire \top_I.branch[5].l_um_iw[246] ;
 wire \top_I.branch[5].l_um_iw[247] ;
 wire \top_I.branch[5].l_um_iw[248] ;
 wire \top_I.branch[5].l_um_iw[249] ;
 wire \top_I.branch[5].l_um_iw[24] ;
 wire \top_I.branch[5].l_um_iw[250] ;
 wire \top_I.branch[5].l_um_iw[251] ;
 wire \top_I.branch[5].l_um_iw[252] ;
 wire \top_I.branch[5].l_um_iw[253] ;
 wire \top_I.branch[5].l_um_iw[254] ;
 wire \top_I.branch[5].l_um_iw[255] ;
 wire \top_I.branch[5].l_um_iw[256] ;
 wire \top_I.branch[5].l_um_iw[257] ;
 wire \top_I.branch[5].l_um_iw[258] ;
 wire \top_I.branch[5].l_um_iw[259] ;
 wire \top_I.branch[5].l_um_iw[25] ;
 wire \top_I.branch[5].l_um_iw[260] ;
 wire \top_I.branch[5].l_um_iw[261] ;
 wire \top_I.branch[5].l_um_iw[262] ;
 wire \top_I.branch[5].l_um_iw[263] ;
 wire \top_I.branch[5].l_um_iw[264] ;
 wire \top_I.branch[5].l_um_iw[265] ;
 wire \top_I.branch[5].l_um_iw[266] ;
 wire \top_I.branch[5].l_um_iw[267] ;
 wire \top_I.branch[5].l_um_iw[268] ;
 wire \top_I.branch[5].l_um_iw[269] ;
 wire \top_I.branch[5].l_um_iw[26] ;
 wire \top_I.branch[5].l_um_iw[270] ;
 wire \top_I.branch[5].l_um_iw[271] ;
 wire \top_I.branch[5].l_um_iw[272] ;
 wire \top_I.branch[5].l_um_iw[273] ;
 wire \top_I.branch[5].l_um_iw[274] ;
 wire \top_I.branch[5].l_um_iw[275] ;
 wire \top_I.branch[5].l_um_iw[276] ;
 wire \top_I.branch[5].l_um_iw[277] ;
 wire \top_I.branch[5].l_um_iw[278] ;
 wire \top_I.branch[5].l_um_iw[279] ;
 wire \top_I.branch[5].l_um_iw[27] ;
 wire \top_I.branch[5].l_um_iw[280] ;
 wire \top_I.branch[5].l_um_iw[281] ;
 wire \top_I.branch[5].l_um_iw[282] ;
 wire \top_I.branch[5].l_um_iw[283] ;
 wire \top_I.branch[5].l_um_iw[284] ;
 wire \top_I.branch[5].l_um_iw[285] ;
 wire \top_I.branch[5].l_um_iw[286] ;
 wire \top_I.branch[5].l_um_iw[287] ;
 wire \top_I.branch[5].l_um_iw[28] ;
 wire \top_I.branch[5].l_um_iw[29] ;
 wire \top_I.branch[5].l_um_iw[2] ;
 wire \top_I.branch[5].l_um_iw[30] ;
 wire \top_I.branch[5].l_um_iw[31] ;
 wire \top_I.branch[5].l_um_iw[32] ;
 wire \top_I.branch[5].l_um_iw[33] ;
 wire \top_I.branch[5].l_um_iw[34] ;
 wire \top_I.branch[5].l_um_iw[35] ;
 wire \top_I.branch[5].l_um_iw[36] ;
 wire \top_I.branch[5].l_um_iw[37] ;
 wire \top_I.branch[5].l_um_iw[38] ;
 wire \top_I.branch[5].l_um_iw[39] ;
 wire \top_I.branch[5].l_um_iw[3] ;
 wire \top_I.branch[5].l_um_iw[40] ;
 wire \top_I.branch[5].l_um_iw[41] ;
 wire \top_I.branch[5].l_um_iw[42] ;
 wire \top_I.branch[5].l_um_iw[43] ;
 wire \top_I.branch[5].l_um_iw[44] ;
 wire \top_I.branch[5].l_um_iw[45] ;
 wire \top_I.branch[5].l_um_iw[46] ;
 wire \top_I.branch[5].l_um_iw[47] ;
 wire \top_I.branch[5].l_um_iw[48] ;
 wire \top_I.branch[5].l_um_iw[49] ;
 wire \top_I.branch[5].l_um_iw[4] ;
 wire \top_I.branch[5].l_um_iw[50] ;
 wire \top_I.branch[5].l_um_iw[51] ;
 wire \top_I.branch[5].l_um_iw[52] ;
 wire \top_I.branch[5].l_um_iw[53] ;
 wire \top_I.branch[5].l_um_iw[54] ;
 wire \top_I.branch[5].l_um_iw[55] ;
 wire \top_I.branch[5].l_um_iw[56] ;
 wire \top_I.branch[5].l_um_iw[57] ;
 wire \top_I.branch[5].l_um_iw[58] ;
 wire \top_I.branch[5].l_um_iw[59] ;
 wire \top_I.branch[5].l_um_iw[5] ;
 wire \top_I.branch[5].l_um_iw[60] ;
 wire \top_I.branch[5].l_um_iw[61] ;
 wire \top_I.branch[5].l_um_iw[62] ;
 wire \top_I.branch[5].l_um_iw[63] ;
 wire \top_I.branch[5].l_um_iw[64] ;
 wire \top_I.branch[5].l_um_iw[65] ;
 wire \top_I.branch[5].l_um_iw[66] ;
 wire \top_I.branch[5].l_um_iw[67] ;
 wire \top_I.branch[5].l_um_iw[68] ;
 wire \top_I.branch[5].l_um_iw[69] ;
 wire \top_I.branch[5].l_um_iw[6] ;
 wire \top_I.branch[5].l_um_iw[70] ;
 wire \top_I.branch[5].l_um_iw[71] ;
 wire \top_I.branch[5].l_um_iw[72] ;
 wire \top_I.branch[5].l_um_iw[73] ;
 wire \top_I.branch[5].l_um_iw[74] ;
 wire \top_I.branch[5].l_um_iw[75] ;
 wire \top_I.branch[5].l_um_iw[76] ;
 wire \top_I.branch[5].l_um_iw[77] ;
 wire \top_I.branch[5].l_um_iw[78] ;
 wire \top_I.branch[5].l_um_iw[79] ;
 wire \top_I.branch[5].l_um_iw[7] ;
 wire \top_I.branch[5].l_um_iw[80] ;
 wire \top_I.branch[5].l_um_iw[81] ;
 wire \top_I.branch[5].l_um_iw[82] ;
 wire \top_I.branch[5].l_um_iw[83] ;
 wire \top_I.branch[5].l_um_iw[84] ;
 wire \top_I.branch[5].l_um_iw[85] ;
 wire \top_I.branch[5].l_um_iw[86] ;
 wire \top_I.branch[5].l_um_iw[87] ;
 wire \top_I.branch[5].l_um_iw[88] ;
 wire \top_I.branch[5].l_um_iw[89] ;
 wire \top_I.branch[5].l_um_iw[8] ;
 wire \top_I.branch[5].l_um_iw[90] ;
 wire \top_I.branch[5].l_um_iw[91] ;
 wire \top_I.branch[5].l_um_iw[92] ;
 wire \top_I.branch[5].l_um_iw[93] ;
 wire \top_I.branch[5].l_um_iw[94] ;
 wire \top_I.branch[5].l_um_iw[95] ;
 wire \top_I.branch[5].l_um_iw[96] ;
 wire \top_I.branch[5].l_um_iw[97] ;
 wire \top_I.branch[5].l_um_iw[98] ;
 wire \top_I.branch[5].l_um_iw[99] ;
 wire \top_I.branch[5].l_um_iw[9] ;
 wire \top_I.branch[5].l_um_k_zero[0] ;
 wire \top_I.branch[5].l_um_k_zero[10] ;
 wire \top_I.branch[5].l_um_k_zero[11] ;
 wire \top_I.branch[5].l_um_k_zero[12] ;
 wire \top_I.branch[5].l_um_k_zero[13] ;
 wire \top_I.branch[5].l_um_k_zero[14] ;
 wire \top_I.branch[5].l_um_k_zero[15] ;
 wire \top_I.branch[5].l_um_k_zero[1] ;
 wire \top_I.branch[5].l_um_k_zero[2] ;
 wire \top_I.branch[5].l_um_k_zero[3] ;
 wire \top_I.branch[5].l_um_k_zero[4] ;
 wire \top_I.branch[5].l_um_k_zero[5] ;
 wire \top_I.branch[5].l_um_k_zero[6] ;
 wire \top_I.branch[5].l_um_k_zero[7] ;
 wire \top_I.branch[5].l_um_k_zero[8] ;
 wire \top_I.branch[5].l_um_k_zero[9] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[6].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[6].l_k_one ;
 wire \top_I.branch[6].l_k_zero ;
 wire \top_I.branch[6].l_um_ena[0] ;
 wire \top_I.branch[6].l_um_ena[10] ;
 wire \top_I.branch[6].l_um_ena[11] ;
 wire \top_I.branch[6].l_um_ena[12] ;
 wire \top_I.branch[6].l_um_ena[13] ;
 wire \top_I.branch[6].l_um_ena[14] ;
 wire \top_I.branch[6].l_um_ena[15] ;
 wire \top_I.branch[6].l_um_ena[1] ;
 wire \top_I.branch[6].l_um_ena[2] ;
 wire \top_I.branch[6].l_um_ena[3] ;
 wire \top_I.branch[6].l_um_ena[4] ;
 wire \top_I.branch[6].l_um_ena[5] ;
 wire \top_I.branch[6].l_um_ena[6] ;
 wire \top_I.branch[6].l_um_ena[7] ;
 wire \top_I.branch[6].l_um_ena[8] ;
 wire \top_I.branch[6].l_um_ena[9] ;
 wire \top_I.branch[6].l_um_iw[0] ;
 wire \top_I.branch[6].l_um_iw[100] ;
 wire \top_I.branch[6].l_um_iw[101] ;
 wire \top_I.branch[6].l_um_iw[102] ;
 wire \top_I.branch[6].l_um_iw[103] ;
 wire \top_I.branch[6].l_um_iw[104] ;
 wire \top_I.branch[6].l_um_iw[105] ;
 wire \top_I.branch[6].l_um_iw[106] ;
 wire \top_I.branch[6].l_um_iw[107] ;
 wire \top_I.branch[6].l_um_iw[108] ;
 wire \top_I.branch[6].l_um_iw[109] ;
 wire \top_I.branch[6].l_um_iw[10] ;
 wire \top_I.branch[6].l_um_iw[110] ;
 wire \top_I.branch[6].l_um_iw[111] ;
 wire \top_I.branch[6].l_um_iw[112] ;
 wire \top_I.branch[6].l_um_iw[113] ;
 wire \top_I.branch[6].l_um_iw[114] ;
 wire \top_I.branch[6].l_um_iw[115] ;
 wire \top_I.branch[6].l_um_iw[116] ;
 wire \top_I.branch[6].l_um_iw[117] ;
 wire \top_I.branch[6].l_um_iw[118] ;
 wire \top_I.branch[6].l_um_iw[119] ;
 wire \top_I.branch[6].l_um_iw[11] ;
 wire \top_I.branch[6].l_um_iw[120] ;
 wire \top_I.branch[6].l_um_iw[121] ;
 wire \top_I.branch[6].l_um_iw[122] ;
 wire \top_I.branch[6].l_um_iw[123] ;
 wire \top_I.branch[6].l_um_iw[124] ;
 wire \top_I.branch[6].l_um_iw[125] ;
 wire \top_I.branch[6].l_um_iw[126] ;
 wire \top_I.branch[6].l_um_iw[127] ;
 wire \top_I.branch[6].l_um_iw[128] ;
 wire \top_I.branch[6].l_um_iw[129] ;
 wire \top_I.branch[6].l_um_iw[12] ;
 wire \top_I.branch[6].l_um_iw[130] ;
 wire \top_I.branch[6].l_um_iw[131] ;
 wire \top_I.branch[6].l_um_iw[132] ;
 wire \top_I.branch[6].l_um_iw[133] ;
 wire \top_I.branch[6].l_um_iw[134] ;
 wire \top_I.branch[6].l_um_iw[135] ;
 wire \top_I.branch[6].l_um_iw[136] ;
 wire \top_I.branch[6].l_um_iw[137] ;
 wire \top_I.branch[6].l_um_iw[138] ;
 wire \top_I.branch[6].l_um_iw[139] ;
 wire \top_I.branch[6].l_um_iw[13] ;
 wire \top_I.branch[6].l_um_iw[140] ;
 wire \top_I.branch[6].l_um_iw[141] ;
 wire \top_I.branch[6].l_um_iw[142] ;
 wire \top_I.branch[6].l_um_iw[143] ;
 wire \top_I.branch[6].l_um_iw[144] ;
 wire \top_I.branch[6].l_um_iw[145] ;
 wire \top_I.branch[6].l_um_iw[146] ;
 wire \top_I.branch[6].l_um_iw[147] ;
 wire \top_I.branch[6].l_um_iw[148] ;
 wire \top_I.branch[6].l_um_iw[149] ;
 wire \top_I.branch[6].l_um_iw[14] ;
 wire \top_I.branch[6].l_um_iw[150] ;
 wire \top_I.branch[6].l_um_iw[151] ;
 wire \top_I.branch[6].l_um_iw[152] ;
 wire \top_I.branch[6].l_um_iw[153] ;
 wire \top_I.branch[6].l_um_iw[154] ;
 wire \top_I.branch[6].l_um_iw[155] ;
 wire \top_I.branch[6].l_um_iw[156] ;
 wire \top_I.branch[6].l_um_iw[157] ;
 wire \top_I.branch[6].l_um_iw[158] ;
 wire \top_I.branch[6].l_um_iw[159] ;
 wire \top_I.branch[6].l_um_iw[15] ;
 wire \top_I.branch[6].l_um_iw[160] ;
 wire \top_I.branch[6].l_um_iw[161] ;
 wire \top_I.branch[6].l_um_iw[162] ;
 wire \top_I.branch[6].l_um_iw[163] ;
 wire \top_I.branch[6].l_um_iw[164] ;
 wire \top_I.branch[6].l_um_iw[165] ;
 wire \top_I.branch[6].l_um_iw[166] ;
 wire \top_I.branch[6].l_um_iw[167] ;
 wire \top_I.branch[6].l_um_iw[168] ;
 wire \top_I.branch[6].l_um_iw[169] ;
 wire \top_I.branch[6].l_um_iw[16] ;
 wire \top_I.branch[6].l_um_iw[170] ;
 wire \top_I.branch[6].l_um_iw[171] ;
 wire \top_I.branch[6].l_um_iw[172] ;
 wire \top_I.branch[6].l_um_iw[173] ;
 wire \top_I.branch[6].l_um_iw[174] ;
 wire \top_I.branch[6].l_um_iw[175] ;
 wire \top_I.branch[6].l_um_iw[176] ;
 wire \top_I.branch[6].l_um_iw[177] ;
 wire \top_I.branch[6].l_um_iw[178] ;
 wire \top_I.branch[6].l_um_iw[179] ;
 wire \top_I.branch[6].l_um_iw[17] ;
 wire \top_I.branch[6].l_um_iw[180] ;
 wire \top_I.branch[6].l_um_iw[181] ;
 wire \top_I.branch[6].l_um_iw[182] ;
 wire \top_I.branch[6].l_um_iw[183] ;
 wire \top_I.branch[6].l_um_iw[184] ;
 wire \top_I.branch[6].l_um_iw[185] ;
 wire \top_I.branch[6].l_um_iw[186] ;
 wire \top_I.branch[6].l_um_iw[187] ;
 wire \top_I.branch[6].l_um_iw[188] ;
 wire \top_I.branch[6].l_um_iw[189] ;
 wire \top_I.branch[6].l_um_iw[18] ;
 wire \top_I.branch[6].l_um_iw[190] ;
 wire \top_I.branch[6].l_um_iw[191] ;
 wire \top_I.branch[6].l_um_iw[192] ;
 wire \top_I.branch[6].l_um_iw[193] ;
 wire \top_I.branch[6].l_um_iw[194] ;
 wire \top_I.branch[6].l_um_iw[195] ;
 wire \top_I.branch[6].l_um_iw[196] ;
 wire \top_I.branch[6].l_um_iw[197] ;
 wire \top_I.branch[6].l_um_iw[198] ;
 wire \top_I.branch[6].l_um_iw[199] ;
 wire \top_I.branch[6].l_um_iw[19] ;
 wire \top_I.branch[6].l_um_iw[1] ;
 wire \top_I.branch[6].l_um_iw[200] ;
 wire \top_I.branch[6].l_um_iw[201] ;
 wire \top_I.branch[6].l_um_iw[202] ;
 wire \top_I.branch[6].l_um_iw[203] ;
 wire \top_I.branch[6].l_um_iw[204] ;
 wire \top_I.branch[6].l_um_iw[205] ;
 wire \top_I.branch[6].l_um_iw[206] ;
 wire \top_I.branch[6].l_um_iw[207] ;
 wire \top_I.branch[6].l_um_iw[208] ;
 wire \top_I.branch[6].l_um_iw[209] ;
 wire \top_I.branch[6].l_um_iw[20] ;
 wire \top_I.branch[6].l_um_iw[210] ;
 wire \top_I.branch[6].l_um_iw[211] ;
 wire \top_I.branch[6].l_um_iw[212] ;
 wire \top_I.branch[6].l_um_iw[213] ;
 wire \top_I.branch[6].l_um_iw[214] ;
 wire \top_I.branch[6].l_um_iw[215] ;
 wire \top_I.branch[6].l_um_iw[216] ;
 wire \top_I.branch[6].l_um_iw[217] ;
 wire \top_I.branch[6].l_um_iw[218] ;
 wire \top_I.branch[6].l_um_iw[219] ;
 wire \top_I.branch[6].l_um_iw[21] ;
 wire \top_I.branch[6].l_um_iw[220] ;
 wire \top_I.branch[6].l_um_iw[221] ;
 wire \top_I.branch[6].l_um_iw[222] ;
 wire \top_I.branch[6].l_um_iw[223] ;
 wire \top_I.branch[6].l_um_iw[224] ;
 wire \top_I.branch[6].l_um_iw[225] ;
 wire \top_I.branch[6].l_um_iw[226] ;
 wire \top_I.branch[6].l_um_iw[227] ;
 wire \top_I.branch[6].l_um_iw[228] ;
 wire \top_I.branch[6].l_um_iw[229] ;
 wire \top_I.branch[6].l_um_iw[22] ;
 wire \top_I.branch[6].l_um_iw[230] ;
 wire \top_I.branch[6].l_um_iw[231] ;
 wire \top_I.branch[6].l_um_iw[232] ;
 wire \top_I.branch[6].l_um_iw[233] ;
 wire \top_I.branch[6].l_um_iw[234] ;
 wire \top_I.branch[6].l_um_iw[235] ;
 wire \top_I.branch[6].l_um_iw[236] ;
 wire \top_I.branch[6].l_um_iw[237] ;
 wire \top_I.branch[6].l_um_iw[238] ;
 wire \top_I.branch[6].l_um_iw[239] ;
 wire \top_I.branch[6].l_um_iw[23] ;
 wire \top_I.branch[6].l_um_iw[240] ;
 wire \top_I.branch[6].l_um_iw[241] ;
 wire \top_I.branch[6].l_um_iw[242] ;
 wire \top_I.branch[6].l_um_iw[243] ;
 wire \top_I.branch[6].l_um_iw[244] ;
 wire \top_I.branch[6].l_um_iw[245] ;
 wire \top_I.branch[6].l_um_iw[246] ;
 wire \top_I.branch[6].l_um_iw[247] ;
 wire \top_I.branch[6].l_um_iw[248] ;
 wire \top_I.branch[6].l_um_iw[249] ;
 wire \top_I.branch[6].l_um_iw[24] ;
 wire \top_I.branch[6].l_um_iw[250] ;
 wire \top_I.branch[6].l_um_iw[251] ;
 wire \top_I.branch[6].l_um_iw[252] ;
 wire \top_I.branch[6].l_um_iw[253] ;
 wire \top_I.branch[6].l_um_iw[254] ;
 wire \top_I.branch[6].l_um_iw[255] ;
 wire \top_I.branch[6].l_um_iw[256] ;
 wire \top_I.branch[6].l_um_iw[257] ;
 wire \top_I.branch[6].l_um_iw[258] ;
 wire \top_I.branch[6].l_um_iw[259] ;
 wire \top_I.branch[6].l_um_iw[25] ;
 wire \top_I.branch[6].l_um_iw[260] ;
 wire \top_I.branch[6].l_um_iw[261] ;
 wire \top_I.branch[6].l_um_iw[262] ;
 wire \top_I.branch[6].l_um_iw[263] ;
 wire \top_I.branch[6].l_um_iw[264] ;
 wire \top_I.branch[6].l_um_iw[265] ;
 wire \top_I.branch[6].l_um_iw[266] ;
 wire \top_I.branch[6].l_um_iw[267] ;
 wire \top_I.branch[6].l_um_iw[268] ;
 wire \top_I.branch[6].l_um_iw[269] ;
 wire \top_I.branch[6].l_um_iw[26] ;
 wire \top_I.branch[6].l_um_iw[270] ;
 wire \top_I.branch[6].l_um_iw[271] ;
 wire \top_I.branch[6].l_um_iw[272] ;
 wire \top_I.branch[6].l_um_iw[273] ;
 wire \top_I.branch[6].l_um_iw[274] ;
 wire \top_I.branch[6].l_um_iw[275] ;
 wire \top_I.branch[6].l_um_iw[276] ;
 wire \top_I.branch[6].l_um_iw[277] ;
 wire \top_I.branch[6].l_um_iw[278] ;
 wire \top_I.branch[6].l_um_iw[279] ;
 wire \top_I.branch[6].l_um_iw[27] ;
 wire \top_I.branch[6].l_um_iw[280] ;
 wire \top_I.branch[6].l_um_iw[281] ;
 wire \top_I.branch[6].l_um_iw[282] ;
 wire \top_I.branch[6].l_um_iw[283] ;
 wire \top_I.branch[6].l_um_iw[284] ;
 wire \top_I.branch[6].l_um_iw[285] ;
 wire \top_I.branch[6].l_um_iw[286] ;
 wire \top_I.branch[6].l_um_iw[287] ;
 wire \top_I.branch[6].l_um_iw[28] ;
 wire \top_I.branch[6].l_um_iw[29] ;
 wire \top_I.branch[6].l_um_iw[2] ;
 wire \top_I.branch[6].l_um_iw[30] ;
 wire \top_I.branch[6].l_um_iw[31] ;
 wire \top_I.branch[6].l_um_iw[32] ;
 wire \top_I.branch[6].l_um_iw[33] ;
 wire \top_I.branch[6].l_um_iw[34] ;
 wire \top_I.branch[6].l_um_iw[35] ;
 wire \top_I.branch[6].l_um_iw[36] ;
 wire \top_I.branch[6].l_um_iw[37] ;
 wire \top_I.branch[6].l_um_iw[38] ;
 wire \top_I.branch[6].l_um_iw[39] ;
 wire \top_I.branch[6].l_um_iw[3] ;
 wire \top_I.branch[6].l_um_iw[40] ;
 wire \top_I.branch[6].l_um_iw[41] ;
 wire \top_I.branch[6].l_um_iw[42] ;
 wire \top_I.branch[6].l_um_iw[43] ;
 wire \top_I.branch[6].l_um_iw[44] ;
 wire \top_I.branch[6].l_um_iw[45] ;
 wire \top_I.branch[6].l_um_iw[46] ;
 wire \top_I.branch[6].l_um_iw[47] ;
 wire \top_I.branch[6].l_um_iw[48] ;
 wire \top_I.branch[6].l_um_iw[49] ;
 wire \top_I.branch[6].l_um_iw[4] ;
 wire \top_I.branch[6].l_um_iw[50] ;
 wire \top_I.branch[6].l_um_iw[51] ;
 wire \top_I.branch[6].l_um_iw[52] ;
 wire \top_I.branch[6].l_um_iw[53] ;
 wire \top_I.branch[6].l_um_iw[54] ;
 wire \top_I.branch[6].l_um_iw[55] ;
 wire \top_I.branch[6].l_um_iw[56] ;
 wire \top_I.branch[6].l_um_iw[57] ;
 wire \top_I.branch[6].l_um_iw[58] ;
 wire \top_I.branch[6].l_um_iw[59] ;
 wire \top_I.branch[6].l_um_iw[5] ;
 wire \top_I.branch[6].l_um_iw[60] ;
 wire \top_I.branch[6].l_um_iw[61] ;
 wire \top_I.branch[6].l_um_iw[62] ;
 wire \top_I.branch[6].l_um_iw[63] ;
 wire \top_I.branch[6].l_um_iw[64] ;
 wire \top_I.branch[6].l_um_iw[65] ;
 wire \top_I.branch[6].l_um_iw[66] ;
 wire \top_I.branch[6].l_um_iw[67] ;
 wire \top_I.branch[6].l_um_iw[68] ;
 wire \top_I.branch[6].l_um_iw[69] ;
 wire \top_I.branch[6].l_um_iw[6] ;
 wire \top_I.branch[6].l_um_iw[70] ;
 wire \top_I.branch[6].l_um_iw[71] ;
 wire \top_I.branch[6].l_um_iw[72] ;
 wire \top_I.branch[6].l_um_iw[73] ;
 wire \top_I.branch[6].l_um_iw[74] ;
 wire \top_I.branch[6].l_um_iw[75] ;
 wire \top_I.branch[6].l_um_iw[76] ;
 wire \top_I.branch[6].l_um_iw[77] ;
 wire \top_I.branch[6].l_um_iw[78] ;
 wire \top_I.branch[6].l_um_iw[79] ;
 wire \top_I.branch[6].l_um_iw[7] ;
 wire \top_I.branch[6].l_um_iw[80] ;
 wire \top_I.branch[6].l_um_iw[81] ;
 wire \top_I.branch[6].l_um_iw[82] ;
 wire \top_I.branch[6].l_um_iw[83] ;
 wire \top_I.branch[6].l_um_iw[84] ;
 wire \top_I.branch[6].l_um_iw[85] ;
 wire \top_I.branch[6].l_um_iw[86] ;
 wire \top_I.branch[6].l_um_iw[87] ;
 wire \top_I.branch[6].l_um_iw[88] ;
 wire \top_I.branch[6].l_um_iw[89] ;
 wire \top_I.branch[6].l_um_iw[8] ;
 wire \top_I.branch[6].l_um_iw[90] ;
 wire \top_I.branch[6].l_um_iw[91] ;
 wire \top_I.branch[6].l_um_iw[92] ;
 wire \top_I.branch[6].l_um_iw[93] ;
 wire \top_I.branch[6].l_um_iw[94] ;
 wire \top_I.branch[6].l_um_iw[95] ;
 wire \top_I.branch[6].l_um_iw[96] ;
 wire \top_I.branch[6].l_um_iw[97] ;
 wire \top_I.branch[6].l_um_iw[98] ;
 wire \top_I.branch[6].l_um_iw[99] ;
 wire \top_I.branch[6].l_um_iw[9] ;
 wire \top_I.branch[6].l_um_k_zero[0] ;
 wire \top_I.branch[6].l_um_k_zero[10] ;
 wire \top_I.branch[6].l_um_k_zero[11] ;
 wire \top_I.branch[6].l_um_k_zero[12] ;
 wire \top_I.branch[6].l_um_k_zero[13] ;
 wire \top_I.branch[6].l_um_k_zero[14] ;
 wire \top_I.branch[6].l_um_k_zero[15] ;
 wire \top_I.branch[6].l_um_k_zero[1] ;
 wire \top_I.branch[6].l_um_k_zero[2] ;
 wire \top_I.branch[6].l_um_k_zero[3] ;
 wire \top_I.branch[6].l_um_k_zero[4] ;
 wire \top_I.branch[6].l_um_k_zero[5] ;
 wire \top_I.branch[6].l_um_k_zero[6] ;
 wire \top_I.branch[6].l_um_k_zero[7] ;
 wire \top_I.branch[6].l_um_k_zero[8] ;
 wire \top_I.branch[6].l_um_k_zero[9] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[0] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[1] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[2] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[3] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[4] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[5] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[6] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_oe[7] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[0] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[1] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[2] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[3] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[4] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[5] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[6] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uio_out[7] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[0] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[1] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[2] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[3] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[4] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[5] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[6] ;
 wire \top_I.branch[7].col_um[0].um_top_I.uo_out[7] ;
 wire \top_I.branch[7].l_k_one ;
 wire \top_I.branch[7].l_k_zero ;
 wire \top_I.branch[7].l_um_ena[0] ;
 wire \top_I.branch[7].l_um_ena[10] ;
 wire \top_I.branch[7].l_um_ena[11] ;
 wire \top_I.branch[7].l_um_ena[12] ;
 wire \top_I.branch[7].l_um_ena[13] ;
 wire \top_I.branch[7].l_um_ena[14] ;
 wire \top_I.branch[7].l_um_ena[15] ;
 wire \top_I.branch[7].l_um_ena[1] ;
 wire \top_I.branch[7].l_um_ena[2] ;
 wire \top_I.branch[7].l_um_ena[3] ;
 wire \top_I.branch[7].l_um_ena[4] ;
 wire \top_I.branch[7].l_um_ena[5] ;
 wire \top_I.branch[7].l_um_ena[6] ;
 wire \top_I.branch[7].l_um_ena[7] ;
 wire \top_I.branch[7].l_um_ena[8] ;
 wire \top_I.branch[7].l_um_ena[9] ;
 wire \top_I.branch[7].l_um_iw[0] ;
 wire \top_I.branch[7].l_um_iw[100] ;
 wire \top_I.branch[7].l_um_iw[101] ;
 wire \top_I.branch[7].l_um_iw[102] ;
 wire \top_I.branch[7].l_um_iw[103] ;
 wire \top_I.branch[7].l_um_iw[104] ;
 wire \top_I.branch[7].l_um_iw[105] ;
 wire \top_I.branch[7].l_um_iw[106] ;
 wire \top_I.branch[7].l_um_iw[107] ;
 wire \top_I.branch[7].l_um_iw[108] ;
 wire \top_I.branch[7].l_um_iw[109] ;
 wire \top_I.branch[7].l_um_iw[10] ;
 wire \top_I.branch[7].l_um_iw[110] ;
 wire \top_I.branch[7].l_um_iw[111] ;
 wire \top_I.branch[7].l_um_iw[112] ;
 wire \top_I.branch[7].l_um_iw[113] ;
 wire \top_I.branch[7].l_um_iw[114] ;
 wire \top_I.branch[7].l_um_iw[115] ;
 wire \top_I.branch[7].l_um_iw[116] ;
 wire \top_I.branch[7].l_um_iw[117] ;
 wire \top_I.branch[7].l_um_iw[118] ;
 wire \top_I.branch[7].l_um_iw[119] ;
 wire \top_I.branch[7].l_um_iw[11] ;
 wire \top_I.branch[7].l_um_iw[120] ;
 wire \top_I.branch[7].l_um_iw[121] ;
 wire \top_I.branch[7].l_um_iw[122] ;
 wire \top_I.branch[7].l_um_iw[123] ;
 wire \top_I.branch[7].l_um_iw[124] ;
 wire \top_I.branch[7].l_um_iw[125] ;
 wire \top_I.branch[7].l_um_iw[126] ;
 wire \top_I.branch[7].l_um_iw[127] ;
 wire \top_I.branch[7].l_um_iw[128] ;
 wire \top_I.branch[7].l_um_iw[129] ;
 wire \top_I.branch[7].l_um_iw[12] ;
 wire \top_I.branch[7].l_um_iw[130] ;
 wire \top_I.branch[7].l_um_iw[131] ;
 wire \top_I.branch[7].l_um_iw[132] ;
 wire \top_I.branch[7].l_um_iw[133] ;
 wire \top_I.branch[7].l_um_iw[134] ;
 wire \top_I.branch[7].l_um_iw[135] ;
 wire \top_I.branch[7].l_um_iw[136] ;
 wire \top_I.branch[7].l_um_iw[137] ;
 wire \top_I.branch[7].l_um_iw[138] ;
 wire \top_I.branch[7].l_um_iw[139] ;
 wire \top_I.branch[7].l_um_iw[13] ;
 wire \top_I.branch[7].l_um_iw[140] ;
 wire \top_I.branch[7].l_um_iw[141] ;
 wire \top_I.branch[7].l_um_iw[142] ;
 wire \top_I.branch[7].l_um_iw[143] ;
 wire \top_I.branch[7].l_um_iw[144] ;
 wire \top_I.branch[7].l_um_iw[145] ;
 wire \top_I.branch[7].l_um_iw[146] ;
 wire \top_I.branch[7].l_um_iw[147] ;
 wire \top_I.branch[7].l_um_iw[148] ;
 wire \top_I.branch[7].l_um_iw[149] ;
 wire \top_I.branch[7].l_um_iw[14] ;
 wire \top_I.branch[7].l_um_iw[150] ;
 wire \top_I.branch[7].l_um_iw[151] ;
 wire \top_I.branch[7].l_um_iw[152] ;
 wire \top_I.branch[7].l_um_iw[153] ;
 wire \top_I.branch[7].l_um_iw[154] ;
 wire \top_I.branch[7].l_um_iw[155] ;
 wire \top_I.branch[7].l_um_iw[156] ;
 wire \top_I.branch[7].l_um_iw[157] ;
 wire \top_I.branch[7].l_um_iw[158] ;
 wire \top_I.branch[7].l_um_iw[159] ;
 wire \top_I.branch[7].l_um_iw[15] ;
 wire \top_I.branch[7].l_um_iw[160] ;
 wire \top_I.branch[7].l_um_iw[161] ;
 wire \top_I.branch[7].l_um_iw[162] ;
 wire \top_I.branch[7].l_um_iw[163] ;
 wire \top_I.branch[7].l_um_iw[164] ;
 wire \top_I.branch[7].l_um_iw[165] ;
 wire \top_I.branch[7].l_um_iw[166] ;
 wire \top_I.branch[7].l_um_iw[167] ;
 wire \top_I.branch[7].l_um_iw[168] ;
 wire \top_I.branch[7].l_um_iw[169] ;
 wire \top_I.branch[7].l_um_iw[16] ;
 wire \top_I.branch[7].l_um_iw[170] ;
 wire \top_I.branch[7].l_um_iw[171] ;
 wire \top_I.branch[7].l_um_iw[172] ;
 wire \top_I.branch[7].l_um_iw[173] ;
 wire \top_I.branch[7].l_um_iw[174] ;
 wire \top_I.branch[7].l_um_iw[175] ;
 wire \top_I.branch[7].l_um_iw[176] ;
 wire \top_I.branch[7].l_um_iw[177] ;
 wire \top_I.branch[7].l_um_iw[178] ;
 wire \top_I.branch[7].l_um_iw[179] ;
 wire \top_I.branch[7].l_um_iw[17] ;
 wire \top_I.branch[7].l_um_iw[180] ;
 wire \top_I.branch[7].l_um_iw[181] ;
 wire \top_I.branch[7].l_um_iw[182] ;
 wire \top_I.branch[7].l_um_iw[183] ;
 wire \top_I.branch[7].l_um_iw[184] ;
 wire \top_I.branch[7].l_um_iw[185] ;
 wire \top_I.branch[7].l_um_iw[186] ;
 wire \top_I.branch[7].l_um_iw[187] ;
 wire \top_I.branch[7].l_um_iw[188] ;
 wire \top_I.branch[7].l_um_iw[189] ;
 wire \top_I.branch[7].l_um_iw[18] ;
 wire \top_I.branch[7].l_um_iw[190] ;
 wire \top_I.branch[7].l_um_iw[191] ;
 wire \top_I.branch[7].l_um_iw[192] ;
 wire \top_I.branch[7].l_um_iw[193] ;
 wire \top_I.branch[7].l_um_iw[194] ;
 wire \top_I.branch[7].l_um_iw[195] ;
 wire \top_I.branch[7].l_um_iw[196] ;
 wire \top_I.branch[7].l_um_iw[197] ;
 wire \top_I.branch[7].l_um_iw[198] ;
 wire \top_I.branch[7].l_um_iw[199] ;
 wire \top_I.branch[7].l_um_iw[19] ;
 wire \top_I.branch[7].l_um_iw[1] ;
 wire \top_I.branch[7].l_um_iw[200] ;
 wire \top_I.branch[7].l_um_iw[201] ;
 wire \top_I.branch[7].l_um_iw[202] ;
 wire \top_I.branch[7].l_um_iw[203] ;
 wire \top_I.branch[7].l_um_iw[204] ;
 wire \top_I.branch[7].l_um_iw[205] ;
 wire \top_I.branch[7].l_um_iw[206] ;
 wire \top_I.branch[7].l_um_iw[207] ;
 wire \top_I.branch[7].l_um_iw[208] ;
 wire \top_I.branch[7].l_um_iw[209] ;
 wire \top_I.branch[7].l_um_iw[20] ;
 wire \top_I.branch[7].l_um_iw[210] ;
 wire \top_I.branch[7].l_um_iw[211] ;
 wire \top_I.branch[7].l_um_iw[212] ;
 wire \top_I.branch[7].l_um_iw[213] ;
 wire \top_I.branch[7].l_um_iw[214] ;
 wire \top_I.branch[7].l_um_iw[215] ;
 wire \top_I.branch[7].l_um_iw[216] ;
 wire \top_I.branch[7].l_um_iw[217] ;
 wire \top_I.branch[7].l_um_iw[218] ;
 wire \top_I.branch[7].l_um_iw[219] ;
 wire \top_I.branch[7].l_um_iw[21] ;
 wire \top_I.branch[7].l_um_iw[220] ;
 wire \top_I.branch[7].l_um_iw[221] ;
 wire \top_I.branch[7].l_um_iw[222] ;
 wire \top_I.branch[7].l_um_iw[223] ;
 wire \top_I.branch[7].l_um_iw[224] ;
 wire \top_I.branch[7].l_um_iw[225] ;
 wire \top_I.branch[7].l_um_iw[226] ;
 wire \top_I.branch[7].l_um_iw[227] ;
 wire \top_I.branch[7].l_um_iw[228] ;
 wire \top_I.branch[7].l_um_iw[229] ;
 wire \top_I.branch[7].l_um_iw[22] ;
 wire \top_I.branch[7].l_um_iw[230] ;
 wire \top_I.branch[7].l_um_iw[231] ;
 wire \top_I.branch[7].l_um_iw[232] ;
 wire \top_I.branch[7].l_um_iw[233] ;
 wire \top_I.branch[7].l_um_iw[234] ;
 wire \top_I.branch[7].l_um_iw[235] ;
 wire \top_I.branch[7].l_um_iw[236] ;
 wire \top_I.branch[7].l_um_iw[237] ;
 wire \top_I.branch[7].l_um_iw[238] ;
 wire \top_I.branch[7].l_um_iw[239] ;
 wire \top_I.branch[7].l_um_iw[23] ;
 wire \top_I.branch[7].l_um_iw[240] ;
 wire \top_I.branch[7].l_um_iw[241] ;
 wire \top_I.branch[7].l_um_iw[242] ;
 wire \top_I.branch[7].l_um_iw[243] ;
 wire \top_I.branch[7].l_um_iw[244] ;
 wire \top_I.branch[7].l_um_iw[245] ;
 wire \top_I.branch[7].l_um_iw[246] ;
 wire \top_I.branch[7].l_um_iw[247] ;
 wire \top_I.branch[7].l_um_iw[248] ;
 wire \top_I.branch[7].l_um_iw[249] ;
 wire \top_I.branch[7].l_um_iw[24] ;
 wire \top_I.branch[7].l_um_iw[250] ;
 wire \top_I.branch[7].l_um_iw[251] ;
 wire \top_I.branch[7].l_um_iw[252] ;
 wire \top_I.branch[7].l_um_iw[253] ;
 wire \top_I.branch[7].l_um_iw[254] ;
 wire \top_I.branch[7].l_um_iw[255] ;
 wire \top_I.branch[7].l_um_iw[256] ;
 wire \top_I.branch[7].l_um_iw[257] ;
 wire \top_I.branch[7].l_um_iw[258] ;
 wire \top_I.branch[7].l_um_iw[259] ;
 wire \top_I.branch[7].l_um_iw[25] ;
 wire \top_I.branch[7].l_um_iw[260] ;
 wire \top_I.branch[7].l_um_iw[261] ;
 wire \top_I.branch[7].l_um_iw[262] ;
 wire \top_I.branch[7].l_um_iw[263] ;
 wire \top_I.branch[7].l_um_iw[264] ;
 wire \top_I.branch[7].l_um_iw[265] ;
 wire \top_I.branch[7].l_um_iw[266] ;
 wire \top_I.branch[7].l_um_iw[267] ;
 wire \top_I.branch[7].l_um_iw[268] ;
 wire \top_I.branch[7].l_um_iw[269] ;
 wire \top_I.branch[7].l_um_iw[26] ;
 wire \top_I.branch[7].l_um_iw[270] ;
 wire \top_I.branch[7].l_um_iw[271] ;
 wire \top_I.branch[7].l_um_iw[272] ;
 wire \top_I.branch[7].l_um_iw[273] ;
 wire \top_I.branch[7].l_um_iw[274] ;
 wire \top_I.branch[7].l_um_iw[275] ;
 wire \top_I.branch[7].l_um_iw[276] ;
 wire \top_I.branch[7].l_um_iw[277] ;
 wire \top_I.branch[7].l_um_iw[278] ;
 wire \top_I.branch[7].l_um_iw[279] ;
 wire \top_I.branch[7].l_um_iw[27] ;
 wire \top_I.branch[7].l_um_iw[280] ;
 wire \top_I.branch[7].l_um_iw[281] ;
 wire \top_I.branch[7].l_um_iw[282] ;
 wire \top_I.branch[7].l_um_iw[283] ;
 wire \top_I.branch[7].l_um_iw[284] ;
 wire \top_I.branch[7].l_um_iw[285] ;
 wire \top_I.branch[7].l_um_iw[286] ;
 wire \top_I.branch[7].l_um_iw[287] ;
 wire \top_I.branch[7].l_um_iw[28] ;
 wire \top_I.branch[7].l_um_iw[29] ;
 wire \top_I.branch[7].l_um_iw[2] ;
 wire \top_I.branch[7].l_um_iw[30] ;
 wire \top_I.branch[7].l_um_iw[31] ;
 wire \top_I.branch[7].l_um_iw[32] ;
 wire \top_I.branch[7].l_um_iw[33] ;
 wire \top_I.branch[7].l_um_iw[34] ;
 wire \top_I.branch[7].l_um_iw[35] ;
 wire \top_I.branch[7].l_um_iw[36] ;
 wire \top_I.branch[7].l_um_iw[37] ;
 wire \top_I.branch[7].l_um_iw[38] ;
 wire \top_I.branch[7].l_um_iw[39] ;
 wire \top_I.branch[7].l_um_iw[3] ;
 wire \top_I.branch[7].l_um_iw[40] ;
 wire \top_I.branch[7].l_um_iw[41] ;
 wire \top_I.branch[7].l_um_iw[42] ;
 wire \top_I.branch[7].l_um_iw[43] ;
 wire \top_I.branch[7].l_um_iw[44] ;
 wire \top_I.branch[7].l_um_iw[45] ;
 wire \top_I.branch[7].l_um_iw[46] ;
 wire \top_I.branch[7].l_um_iw[47] ;
 wire \top_I.branch[7].l_um_iw[48] ;
 wire \top_I.branch[7].l_um_iw[49] ;
 wire \top_I.branch[7].l_um_iw[4] ;
 wire \top_I.branch[7].l_um_iw[50] ;
 wire \top_I.branch[7].l_um_iw[51] ;
 wire \top_I.branch[7].l_um_iw[52] ;
 wire \top_I.branch[7].l_um_iw[53] ;
 wire \top_I.branch[7].l_um_iw[54] ;
 wire \top_I.branch[7].l_um_iw[55] ;
 wire \top_I.branch[7].l_um_iw[56] ;
 wire \top_I.branch[7].l_um_iw[57] ;
 wire \top_I.branch[7].l_um_iw[58] ;
 wire \top_I.branch[7].l_um_iw[59] ;
 wire \top_I.branch[7].l_um_iw[5] ;
 wire \top_I.branch[7].l_um_iw[60] ;
 wire \top_I.branch[7].l_um_iw[61] ;
 wire \top_I.branch[7].l_um_iw[62] ;
 wire \top_I.branch[7].l_um_iw[63] ;
 wire \top_I.branch[7].l_um_iw[64] ;
 wire \top_I.branch[7].l_um_iw[65] ;
 wire \top_I.branch[7].l_um_iw[66] ;
 wire \top_I.branch[7].l_um_iw[67] ;
 wire \top_I.branch[7].l_um_iw[68] ;
 wire \top_I.branch[7].l_um_iw[69] ;
 wire \top_I.branch[7].l_um_iw[6] ;
 wire \top_I.branch[7].l_um_iw[70] ;
 wire \top_I.branch[7].l_um_iw[71] ;
 wire \top_I.branch[7].l_um_iw[72] ;
 wire \top_I.branch[7].l_um_iw[73] ;
 wire \top_I.branch[7].l_um_iw[74] ;
 wire \top_I.branch[7].l_um_iw[75] ;
 wire \top_I.branch[7].l_um_iw[76] ;
 wire \top_I.branch[7].l_um_iw[77] ;
 wire \top_I.branch[7].l_um_iw[78] ;
 wire \top_I.branch[7].l_um_iw[79] ;
 wire \top_I.branch[7].l_um_iw[7] ;
 wire \top_I.branch[7].l_um_iw[80] ;
 wire \top_I.branch[7].l_um_iw[81] ;
 wire \top_I.branch[7].l_um_iw[82] ;
 wire \top_I.branch[7].l_um_iw[83] ;
 wire \top_I.branch[7].l_um_iw[84] ;
 wire \top_I.branch[7].l_um_iw[85] ;
 wire \top_I.branch[7].l_um_iw[86] ;
 wire \top_I.branch[7].l_um_iw[87] ;
 wire \top_I.branch[7].l_um_iw[88] ;
 wire \top_I.branch[7].l_um_iw[89] ;
 wire \top_I.branch[7].l_um_iw[8] ;
 wire \top_I.branch[7].l_um_iw[90] ;
 wire \top_I.branch[7].l_um_iw[91] ;
 wire \top_I.branch[7].l_um_iw[92] ;
 wire \top_I.branch[7].l_um_iw[93] ;
 wire \top_I.branch[7].l_um_iw[94] ;
 wire \top_I.branch[7].l_um_iw[95] ;
 wire \top_I.branch[7].l_um_iw[96] ;
 wire \top_I.branch[7].l_um_iw[97] ;
 wire \top_I.branch[7].l_um_iw[98] ;
 wire \top_I.branch[7].l_um_iw[99] ;
 wire \top_I.branch[7].l_um_iw[9] ;
 wire \top_I.branch[7].l_um_k_zero[0] ;
 wire \top_I.branch[7].l_um_k_zero[10] ;
 wire \top_I.branch[7].l_um_k_zero[11] ;
 wire \top_I.branch[7].l_um_k_zero[12] ;
 wire \top_I.branch[7].l_um_k_zero[13] ;
 wire \top_I.branch[7].l_um_k_zero[14] ;
 wire \top_I.branch[7].l_um_k_zero[15] ;
 wire \top_I.branch[7].l_um_k_zero[1] ;
 wire \top_I.branch[7].l_um_k_zero[2] ;
 wire \top_I.branch[7].l_um_k_zero[3] ;
 wire \top_I.branch[7].l_um_k_zero[4] ;
 wire \top_I.branch[7].l_um_k_zero[5] ;
 wire \top_I.branch[7].l_um_k_zero[6] ;
 wire \top_I.branch[7].l_um_k_zero[7] ;
 wire \top_I.branch[7].l_um_k_zero[8] ;
 wire \top_I.branch[7].l_um_k_zero[9] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[8].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[8].l_k_one ;
 wire \top_I.branch[8].l_k_zero ;
 wire \top_I.branch[8].l_um_ena[0] ;
 wire \top_I.branch[8].l_um_ena[10] ;
 wire \top_I.branch[8].l_um_ena[11] ;
 wire \top_I.branch[8].l_um_ena[12] ;
 wire \top_I.branch[8].l_um_ena[13] ;
 wire \top_I.branch[8].l_um_ena[14] ;
 wire \top_I.branch[8].l_um_ena[15] ;
 wire \top_I.branch[8].l_um_ena[1] ;
 wire \top_I.branch[8].l_um_ena[2] ;
 wire \top_I.branch[8].l_um_ena[3] ;
 wire \top_I.branch[8].l_um_ena[4] ;
 wire \top_I.branch[8].l_um_ena[5] ;
 wire \top_I.branch[8].l_um_ena[6] ;
 wire \top_I.branch[8].l_um_ena[7] ;
 wire \top_I.branch[8].l_um_ena[8] ;
 wire \top_I.branch[8].l_um_ena[9] ;
 wire \top_I.branch[8].l_um_iw[0] ;
 wire \top_I.branch[8].l_um_iw[100] ;
 wire \top_I.branch[8].l_um_iw[101] ;
 wire \top_I.branch[8].l_um_iw[102] ;
 wire \top_I.branch[8].l_um_iw[103] ;
 wire \top_I.branch[8].l_um_iw[104] ;
 wire \top_I.branch[8].l_um_iw[105] ;
 wire \top_I.branch[8].l_um_iw[106] ;
 wire \top_I.branch[8].l_um_iw[107] ;
 wire \top_I.branch[8].l_um_iw[108] ;
 wire \top_I.branch[8].l_um_iw[109] ;
 wire \top_I.branch[8].l_um_iw[10] ;
 wire \top_I.branch[8].l_um_iw[110] ;
 wire \top_I.branch[8].l_um_iw[111] ;
 wire \top_I.branch[8].l_um_iw[112] ;
 wire \top_I.branch[8].l_um_iw[113] ;
 wire \top_I.branch[8].l_um_iw[114] ;
 wire \top_I.branch[8].l_um_iw[115] ;
 wire \top_I.branch[8].l_um_iw[116] ;
 wire \top_I.branch[8].l_um_iw[117] ;
 wire \top_I.branch[8].l_um_iw[118] ;
 wire \top_I.branch[8].l_um_iw[119] ;
 wire \top_I.branch[8].l_um_iw[11] ;
 wire \top_I.branch[8].l_um_iw[120] ;
 wire \top_I.branch[8].l_um_iw[121] ;
 wire \top_I.branch[8].l_um_iw[122] ;
 wire \top_I.branch[8].l_um_iw[123] ;
 wire \top_I.branch[8].l_um_iw[124] ;
 wire \top_I.branch[8].l_um_iw[125] ;
 wire \top_I.branch[8].l_um_iw[126] ;
 wire \top_I.branch[8].l_um_iw[127] ;
 wire \top_I.branch[8].l_um_iw[128] ;
 wire \top_I.branch[8].l_um_iw[129] ;
 wire \top_I.branch[8].l_um_iw[12] ;
 wire \top_I.branch[8].l_um_iw[130] ;
 wire \top_I.branch[8].l_um_iw[131] ;
 wire \top_I.branch[8].l_um_iw[132] ;
 wire \top_I.branch[8].l_um_iw[133] ;
 wire \top_I.branch[8].l_um_iw[134] ;
 wire \top_I.branch[8].l_um_iw[135] ;
 wire \top_I.branch[8].l_um_iw[136] ;
 wire \top_I.branch[8].l_um_iw[137] ;
 wire \top_I.branch[8].l_um_iw[138] ;
 wire \top_I.branch[8].l_um_iw[139] ;
 wire \top_I.branch[8].l_um_iw[13] ;
 wire \top_I.branch[8].l_um_iw[140] ;
 wire \top_I.branch[8].l_um_iw[141] ;
 wire \top_I.branch[8].l_um_iw[142] ;
 wire \top_I.branch[8].l_um_iw[143] ;
 wire \top_I.branch[8].l_um_iw[144] ;
 wire \top_I.branch[8].l_um_iw[145] ;
 wire \top_I.branch[8].l_um_iw[146] ;
 wire \top_I.branch[8].l_um_iw[147] ;
 wire \top_I.branch[8].l_um_iw[148] ;
 wire \top_I.branch[8].l_um_iw[149] ;
 wire \top_I.branch[8].l_um_iw[14] ;
 wire \top_I.branch[8].l_um_iw[150] ;
 wire \top_I.branch[8].l_um_iw[151] ;
 wire \top_I.branch[8].l_um_iw[152] ;
 wire \top_I.branch[8].l_um_iw[153] ;
 wire \top_I.branch[8].l_um_iw[154] ;
 wire \top_I.branch[8].l_um_iw[155] ;
 wire \top_I.branch[8].l_um_iw[156] ;
 wire \top_I.branch[8].l_um_iw[157] ;
 wire \top_I.branch[8].l_um_iw[158] ;
 wire \top_I.branch[8].l_um_iw[159] ;
 wire \top_I.branch[8].l_um_iw[15] ;
 wire \top_I.branch[8].l_um_iw[160] ;
 wire \top_I.branch[8].l_um_iw[161] ;
 wire \top_I.branch[8].l_um_iw[162] ;
 wire \top_I.branch[8].l_um_iw[163] ;
 wire \top_I.branch[8].l_um_iw[164] ;
 wire \top_I.branch[8].l_um_iw[165] ;
 wire \top_I.branch[8].l_um_iw[166] ;
 wire \top_I.branch[8].l_um_iw[167] ;
 wire \top_I.branch[8].l_um_iw[168] ;
 wire \top_I.branch[8].l_um_iw[169] ;
 wire \top_I.branch[8].l_um_iw[16] ;
 wire \top_I.branch[8].l_um_iw[170] ;
 wire \top_I.branch[8].l_um_iw[171] ;
 wire \top_I.branch[8].l_um_iw[172] ;
 wire \top_I.branch[8].l_um_iw[173] ;
 wire \top_I.branch[8].l_um_iw[174] ;
 wire \top_I.branch[8].l_um_iw[175] ;
 wire \top_I.branch[8].l_um_iw[176] ;
 wire \top_I.branch[8].l_um_iw[177] ;
 wire \top_I.branch[8].l_um_iw[178] ;
 wire \top_I.branch[8].l_um_iw[179] ;
 wire \top_I.branch[8].l_um_iw[17] ;
 wire \top_I.branch[8].l_um_iw[180] ;
 wire \top_I.branch[8].l_um_iw[181] ;
 wire \top_I.branch[8].l_um_iw[182] ;
 wire \top_I.branch[8].l_um_iw[183] ;
 wire \top_I.branch[8].l_um_iw[184] ;
 wire \top_I.branch[8].l_um_iw[185] ;
 wire \top_I.branch[8].l_um_iw[186] ;
 wire \top_I.branch[8].l_um_iw[187] ;
 wire \top_I.branch[8].l_um_iw[188] ;
 wire \top_I.branch[8].l_um_iw[189] ;
 wire \top_I.branch[8].l_um_iw[18] ;
 wire \top_I.branch[8].l_um_iw[190] ;
 wire \top_I.branch[8].l_um_iw[191] ;
 wire \top_I.branch[8].l_um_iw[192] ;
 wire \top_I.branch[8].l_um_iw[193] ;
 wire \top_I.branch[8].l_um_iw[194] ;
 wire \top_I.branch[8].l_um_iw[195] ;
 wire \top_I.branch[8].l_um_iw[196] ;
 wire \top_I.branch[8].l_um_iw[197] ;
 wire \top_I.branch[8].l_um_iw[198] ;
 wire \top_I.branch[8].l_um_iw[199] ;
 wire \top_I.branch[8].l_um_iw[19] ;
 wire \top_I.branch[8].l_um_iw[1] ;
 wire \top_I.branch[8].l_um_iw[200] ;
 wire \top_I.branch[8].l_um_iw[201] ;
 wire \top_I.branch[8].l_um_iw[202] ;
 wire \top_I.branch[8].l_um_iw[203] ;
 wire \top_I.branch[8].l_um_iw[204] ;
 wire \top_I.branch[8].l_um_iw[205] ;
 wire \top_I.branch[8].l_um_iw[206] ;
 wire \top_I.branch[8].l_um_iw[207] ;
 wire \top_I.branch[8].l_um_iw[208] ;
 wire \top_I.branch[8].l_um_iw[209] ;
 wire \top_I.branch[8].l_um_iw[20] ;
 wire \top_I.branch[8].l_um_iw[210] ;
 wire \top_I.branch[8].l_um_iw[211] ;
 wire \top_I.branch[8].l_um_iw[212] ;
 wire \top_I.branch[8].l_um_iw[213] ;
 wire \top_I.branch[8].l_um_iw[214] ;
 wire \top_I.branch[8].l_um_iw[215] ;
 wire \top_I.branch[8].l_um_iw[216] ;
 wire \top_I.branch[8].l_um_iw[217] ;
 wire \top_I.branch[8].l_um_iw[218] ;
 wire \top_I.branch[8].l_um_iw[219] ;
 wire \top_I.branch[8].l_um_iw[21] ;
 wire \top_I.branch[8].l_um_iw[220] ;
 wire \top_I.branch[8].l_um_iw[221] ;
 wire \top_I.branch[8].l_um_iw[222] ;
 wire \top_I.branch[8].l_um_iw[223] ;
 wire \top_I.branch[8].l_um_iw[224] ;
 wire \top_I.branch[8].l_um_iw[225] ;
 wire \top_I.branch[8].l_um_iw[226] ;
 wire \top_I.branch[8].l_um_iw[227] ;
 wire \top_I.branch[8].l_um_iw[228] ;
 wire \top_I.branch[8].l_um_iw[229] ;
 wire \top_I.branch[8].l_um_iw[22] ;
 wire \top_I.branch[8].l_um_iw[230] ;
 wire \top_I.branch[8].l_um_iw[231] ;
 wire \top_I.branch[8].l_um_iw[232] ;
 wire \top_I.branch[8].l_um_iw[233] ;
 wire \top_I.branch[8].l_um_iw[234] ;
 wire \top_I.branch[8].l_um_iw[235] ;
 wire \top_I.branch[8].l_um_iw[236] ;
 wire \top_I.branch[8].l_um_iw[237] ;
 wire \top_I.branch[8].l_um_iw[238] ;
 wire \top_I.branch[8].l_um_iw[239] ;
 wire \top_I.branch[8].l_um_iw[23] ;
 wire \top_I.branch[8].l_um_iw[240] ;
 wire \top_I.branch[8].l_um_iw[241] ;
 wire \top_I.branch[8].l_um_iw[242] ;
 wire \top_I.branch[8].l_um_iw[243] ;
 wire \top_I.branch[8].l_um_iw[244] ;
 wire \top_I.branch[8].l_um_iw[245] ;
 wire \top_I.branch[8].l_um_iw[246] ;
 wire \top_I.branch[8].l_um_iw[247] ;
 wire \top_I.branch[8].l_um_iw[248] ;
 wire \top_I.branch[8].l_um_iw[249] ;
 wire \top_I.branch[8].l_um_iw[24] ;
 wire \top_I.branch[8].l_um_iw[250] ;
 wire \top_I.branch[8].l_um_iw[251] ;
 wire \top_I.branch[8].l_um_iw[252] ;
 wire \top_I.branch[8].l_um_iw[253] ;
 wire \top_I.branch[8].l_um_iw[254] ;
 wire \top_I.branch[8].l_um_iw[255] ;
 wire \top_I.branch[8].l_um_iw[256] ;
 wire \top_I.branch[8].l_um_iw[257] ;
 wire \top_I.branch[8].l_um_iw[258] ;
 wire \top_I.branch[8].l_um_iw[259] ;
 wire \top_I.branch[8].l_um_iw[25] ;
 wire \top_I.branch[8].l_um_iw[260] ;
 wire \top_I.branch[8].l_um_iw[261] ;
 wire \top_I.branch[8].l_um_iw[262] ;
 wire \top_I.branch[8].l_um_iw[263] ;
 wire \top_I.branch[8].l_um_iw[264] ;
 wire \top_I.branch[8].l_um_iw[265] ;
 wire \top_I.branch[8].l_um_iw[266] ;
 wire \top_I.branch[8].l_um_iw[267] ;
 wire \top_I.branch[8].l_um_iw[268] ;
 wire \top_I.branch[8].l_um_iw[269] ;
 wire \top_I.branch[8].l_um_iw[26] ;
 wire \top_I.branch[8].l_um_iw[270] ;
 wire \top_I.branch[8].l_um_iw[271] ;
 wire \top_I.branch[8].l_um_iw[272] ;
 wire \top_I.branch[8].l_um_iw[273] ;
 wire \top_I.branch[8].l_um_iw[274] ;
 wire \top_I.branch[8].l_um_iw[275] ;
 wire \top_I.branch[8].l_um_iw[276] ;
 wire \top_I.branch[8].l_um_iw[277] ;
 wire \top_I.branch[8].l_um_iw[278] ;
 wire \top_I.branch[8].l_um_iw[279] ;
 wire \top_I.branch[8].l_um_iw[27] ;
 wire \top_I.branch[8].l_um_iw[280] ;
 wire \top_I.branch[8].l_um_iw[281] ;
 wire \top_I.branch[8].l_um_iw[282] ;
 wire \top_I.branch[8].l_um_iw[283] ;
 wire \top_I.branch[8].l_um_iw[284] ;
 wire \top_I.branch[8].l_um_iw[285] ;
 wire \top_I.branch[8].l_um_iw[286] ;
 wire \top_I.branch[8].l_um_iw[287] ;
 wire \top_I.branch[8].l_um_iw[28] ;
 wire \top_I.branch[8].l_um_iw[29] ;
 wire \top_I.branch[8].l_um_iw[2] ;
 wire \top_I.branch[8].l_um_iw[30] ;
 wire \top_I.branch[8].l_um_iw[31] ;
 wire \top_I.branch[8].l_um_iw[32] ;
 wire \top_I.branch[8].l_um_iw[33] ;
 wire \top_I.branch[8].l_um_iw[34] ;
 wire \top_I.branch[8].l_um_iw[35] ;
 wire \top_I.branch[8].l_um_iw[36] ;
 wire \top_I.branch[8].l_um_iw[37] ;
 wire \top_I.branch[8].l_um_iw[38] ;
 wire \top_I.branch[8].l_um_iw[39] ;
 wire \top_I.branch[8].l_um_iw[3] ;
 wire \top_I.branch[8].l_um_iw[40] ;
 wire \top_I.branch[8].l_um_iw[41] ;
 wire \top_I.branch[8].l_um_iw[42] ;
 wire \top_I.branch[8].l_um_iw[43] ;
 wire \top_I.branch[8].l_um_iw[44] ;
 wire \top_I.branch[8].l_um_iw[45] ;
 wire \top_I.branch[8].l_um_iw[46] ;
 wire \top_I.branch[8].l_um_iw[47] ;
 wire \top_I.branch[8].l_um_iw[48] ;
 wire \top_I.branch[8].l_um_iw[49] ;
 wire \top_I.branch[8].l_um_iw[4] ;
 wire \top_I.branch[8].l_um_iw[50] ;
 wire \top_I.branch[8].l_um_iw[51] ;
 wire \top_I.branch[8].l_um_iw[52] ;
 wire \top_I.branch[8].l_um_iw[53] ;
 wire \top_I.branch[8].l_um_iw[54] ;
 wire \top_I.branch[8].l_um_iw[55] ;
 wire \top_I.branch[8].l_um_iw[56] ;
 wire \top_I.branch[8].l_um_iw[57] ;
 wire \top_I.branch[8].l_um_iw[58] ;
 wire \top_I.branch[8].l_um_iw[59] ;
 wire \top_I.branch[8].l_um_iw[5] ;
 wire \top_I.branch[8].l_um_iw[60] ;
 wire \top_I.branch[8].l_um_iw[61] ;
 wire \top_I.branch[8].l_um_iw[62] ;
 wire \top_I.branch[8].l_um_iw[63] ;
 wire \top_I.branch[8].l_um_iw[64] ;
 wire \top_I.branch[8].l_um_iw[65] ;
 wire \top_I.branch[8].l_um_iw[66] ;
 wire \top_I.branch[8].l_um_iw[67] ;
 wire \top_I.branch[8].l_um_iw[68] ;
 wire \top_I.branch[8].l_um_iw[69] ;
 wire \top_I.branch[8].l_um_iw[6] ;
 wire \top_I.branch[8].l_um_iw[70] ;
 wire \top_I.branch[8].l_um_iw[71] ;
 wire \top_I.branch[8].l_um_iw[72] ;
 wire \top_I.branch[8].l_um_iw[73] ;
 wire \top_I.branch[8].l_um_iw[74] ;
 wire \top_I.branch[8].l_um_iw[75] ;
 wire \top_I.branch[8].l_um_iw[76] ;
 wire \top_I.branch[8].l_um_iw[77] ;
 wire \top_I.branch[8].l_um_iw[78] ;
 wire \top_I.branch[8].l_um_iw[79] ;
 wire \top_I.branch[8].l_um_iw[7] ;
 wire \top_I.branch[8].l_um_iw[80] ;
 wire \top_I.branch[8].l_um_iw[81] ;
 wire \top_I.branch[8].l_um_iw[82] ;
 wire \top_I.branch[8].l_um_iw[83] ;
 wire \top_I.branch[8].l_um_iw[84] ;
 wire \top_I.branch[8].l_um_iw[85] ;
 wire \top_I.branch[8].l_um_iw[86] ;
 wire \top_I.branch[8].l_um_iw[87] ;
 wire \top_I.branch[8].l_um_iw[88] ;
 wire \top_I.branch[8].l_um_iw[89] ;
 wire \top_I.branch[8].l_um_iw[8] ;
 wire \top_I.branch[8].l_um_iw[90] ;
 wire \top_I.branch[8].l_um_iw[91] ;
 wire \top_I.branch[8].l_um_iw[92] ;
 wire \top_I.branch[8].l_um_iw[93] ;
 wire \top_I.branch[8].l_um_iw[94] ;
 wire \top_I.branch[8].l_um_iw[95] ;
 wire \top_I.branch[8].l_um_iw[96] ;
 wire \top_I.branch[8].l_um_iw[97] ;
 wire \top_I.branch[8].l_um_iw[98] ;
 wire \top_I.branch[8].l_um_iw[99] ;
 wire \top_I.branch[8].l_um_iw[9] ;
 wire \top_I.branch[8].l_um_k_zero[0] ;
 wire \top_I.branch[8].l_um_k_zero[10] ;
 wire \top_I.branch[8].l_um_k_zero[11] ;
 wire \top_I.branch[8].l_um_k_zero[12] ;
 wire \top_I.branch[8].l_um_k_zero[13] ;
 wire \top_I.branch[8].l_um_k_zero[14] ;
 wire \top_I.branch[8].l_um_k_zero[15] ;
 wire \top_I.branch[8].l_um_k_zero[1] ;
 wire \top_I.branch[8].l_um_k_zero[2] ;
 wire \top_I.branch[8].l_um_k_zero[3] ;
 wire \top_I.branch[8].l_um_k_zero[4] ;
 wire \top_I.branch[8].l_um_k_zero[5] ;
 wire \top_I.branch[8].l_um_k_zero[6] ;
 wire \top_I.branch[8].l_um_k_zero[7] ;
 wire \top_I.branch[8].l_um_k_zero[8] ;
 wire \top_I.branch[8].l_um_k_zero[9] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[0] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[1] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[2] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[3] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[4] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[5] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[6] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_oe[7] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[0] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[1] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[2] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[3] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[4] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[5] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[6] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uio_out[7] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[0] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[1] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[2] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[3] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[4] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[5] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[6] ;
 wire \top_I.branch[9].col_um[0].um_bot_I.uo_out[7] ;
 wire \top_I.branch[9].l_k_one ;
 wire \top_I.branch[9].l_k_zero ;
 wire \top_I.branch[9].l_um_ena[0] ;
 wire \top_I.branch[9].l_um_ena[10] ;
 wire \top_I.branch[9].l_um_ena[11] ;
 wire \top_I.branch[9].l_um_ena[12] ;
 wire \top_I.branch[9].l_um_ena[13] ;
 wire \top_I.branch[9].l_um_ena[14] ;
 wire \top_I.branch[9].l_um_ena[15] ;
 wire \top_I.branch[9].l_um_ena[1] ;
 wire \top_I.branch[9].l_um_ena[2] ;
 wire \top_I.branch[9].l_um_ena[3] ;
 wire \top_I.branch[9].l_um_ena[4] ;
 wire \top_I.branch[9].l_um_ena[5] ;
 wire \top_I.branch[9].l_um_ena[6] ;
 wire \top_I.branch[9].l_um_ena[7] ;
 wire \top_I.branch[9].l_um_ena[8] ;
 wire \top_I.branch[9].l_um_ena[9] ;
 wire \top_I.branch[9].l_um_iw[0] ;
 wire \top_I.branch[9].l_um_iw[100] ;
 wire \top_I.branch[9].l_um_iw[101] ;
 wire \top_I.branch[9].l_um_iw[102] ;
 wire \top_I.branch[9].l_um_iw[103] ;
 wire \top_I.branch[9].l_um_iw[104] ;
 wire \top_I.branch[9].l_um_iw[105] ;
 wire \top_I.branch[9].l_um_iw[106] ;
 wire \top_I.branch[9].l_um_iw[107] ;
 wire \top_I.branch[9].l_um_iw[108] ;
 wire \top_I.branch[9].l_um_iw[109] ;
 wire \top_I.branch[9].l_um_iw[10] ;
 wire \top_I.branch[9].l_um_iw[110] ;
 wire \top_I.branch[9].l_um_iw[111] ;
 wire \top_I.branch[9].l_um_iw[112] ;
 wire \top_I.branch[9].l_um_iw[113] ;
 wire \top_I.branch[9].l_um_iw[114] ;
 wire \top_I.branch[9].l_um_iw[115] ;
 wire \top_I.branch[9].l_um_iw[116] ;
 wire \top_I.branch[9].l_um_iw[117] ;
 wire \top_I.branch[9].l_um_iw[118] ;
 wire \top_I.branch[9].l_um_iw[119] ;
 wire \top_I.branch[9].l_um_iw[11] ;
 wire \top_I.branch[9].l_um_iw[120] ;
 wire \top_I.branch[9].l_um_iw[121] ;
 wire \top_I.branch[9].l_um_iw[122] ;
 wire \top_I.branch[9].l_um_iw[123] ;
 wire \top_I.branch[9].l_um_iw[124] ;
 wire \top_I.branch[9].l_um_iw[125] ;
 wire \top_I.branch[9].l_um_iw[126] ;
 wire \top_I.branch[9].l_um_iw[127] ;
 wire \top_I.branch[9].l_um_iw[128] ;
 wire \top_I.branch[9].l_um_iw[129] ;
 wire \top_I.branch[9].l_um_iw[12] ;
 wire \top_I.branch[9].l_um_iw[130] ;
 wire \top_I.branch[9].l_um_iw[131] ;
 wire \top_I.branch[9].l_um_iw[132] ;
 wire \top_I.branch[9].l_um_iw[133] ;
 wire \top_I.branch[9].l_um_iw[134] ;
 wire \top_I.branch[9].l_um_iw[135] ;
 wire \top_I.branch[9].l_um_iw[136] ;
 wire \top_I.branch[9].l_um_iw[137] ;
 wire \top_I.branch[9].l_um_iw[138] ;
 wire \top_I.branch[9].l_um_iw[139] ;
 wire \top_I.branch[9].l_um_iw[13] ;
 wire \top_I.branch[9].l_um_iw[140] ;
 wire \top_I.branch[9].l_um_iw[141] ;
 wire \top_I.branch[9].l_um_iw[142] ;
 wire \top_I.branch[9].l_um_iw[143] ;
 wire \top_I.branch[9].l_um_iw[144] ;
 wire \top_I.branch[9].l_um_iw[145] ;
 wire \top_I.branch[9].l_um_iw[146] ;
 wire \top_I.branch[9].l_um_iw[147] ;
 wire \top_I.branch[9].l_um_iw[148] ;
 wire \top_I.branch[9].l_um_iw[149] ;
 wire \top_I.branch[9].l_um_iw[14] ;
 wire \top_I.branch[9].l_um_iw[150] ;
 wire \top_I.branch[9].l_um_iw[151] ;
 wire \top_I.branch[9].l_um_iw[152] ;
 wire \top_I.branch[9].l_um_iw[153] ;
 wire \top_I.branch[9].l_um_iw[154] ;
 wire \top_I.branch[9].l_um_iw[155] ;
 wire \top_I.branch[9].l_um_iw[156] ;
 wire \top_I.branch[9].l_um_iw[157] ;
 wire \top_I.branch[9].l_um_iw[158] ;
 wire \top_I.branch[9].l_um_iw[159] ;
 wire \top_I.branch[9].l_um_iw[15] ;
 wire \top_I.branch[9].l_um_iw[160] ;
 wire \top_I.branch[9].l_um_iw[161] ;
 wire \top_I.branch[9].l_um_iw[162] ;
 wire \top_I.branch[9].l_um_iw[163] ;
 wire \top_I.branch[9].l_um_iw[164] ;
 wire \top_I.branch[9].l_um_iw[165] ;
 wire \top_I.branch[9].l_um_iw[166] ;
 wire \top_I.branch[9].l_um_iw[167] ;
 wire \top_I.branch[9].l_um_iw[168] ;
 wire \top_I.branch[9].l_um_iw[169] ;
 wire \top_I.branch[9].l_um_iw[16] ;
 wire \top_I.branch[9].l_um_iw[170] ;
 wire \top_I.branch[9].l_um_iw[171] ;
 wire \top_I.branch[9].l_um_iw[172] ;
 wire \top_I.branch[9].l_um_iw[173] ;
 wire \top_I.branch[9].l_um_iw[174] ;
 wire \top_I.branch[9].l_um_iw[175] ;
 wire \top_I.branch[9].l_um_iw[176] ;
 wire \top_I.branch[9].l_um_iw[177] ;
 wire \top_I.branch[9].l_um_iw[178] ;
 wire \top_I.branch[9].l_um_iw[179] ;
 wire \top_I.branch[9].l_um_iw[17] ;
 wire \top_I.branch[9].l_um_iw[180] ;
 wire \top_I.branch[9].l_um_iw[181] ;
 wire \top_I.branch[9].l_um_iw[182] ;
 wire \top_I.branch[9].l_um_iw[183] ;
 wire \top_I.branch[9].l_um_iw[184] ;
 wire \top_I.branch[9].l_um_iw[185] ;
 wire \top_I.branch[9].l_um_iw[186] ;
 wire \top_I.branch[9].l_um_iw[187] ;
 wire \top_I.branch[9].l_um_iw[188] ;
 wire \top_I.branch[9].l_um_iw[189] ;
 wire \top_I.branch[9].l_um_iw[18] ;
 wire \top_I.branch[9].l_um_iw[190] ;
 wire \top_I.branch[9].l_um_iw[191] ;
 wire \top_I.branch[9].l_um_iw[192] ;
 wire \top_I.branch[9].l_um_iw[193] ;
 wire \top_I.branch[9].l_um_iw[194] ;
 wire \top_I.branch[9].l_um_iw[195] ;
 wire \top_I.branch[9].l_um_iw[196] ;
 wire \top_I.branch[9].l_um_iw[197] ;
 wire \top_I.branch[9].l_um_iw[198] ;
 wire \top_I.branch[9].l_um_iw[199] ;
 wire \top_I.branch[9].l_um_iw[19] ;
 wire \top_I.branch[9].l_um_iw[1] ;
 wire \top_I.branch[9].l_um_iw[200] ;
 wire \top_I.branch[9].l_um_iw[201] ;
 wire \top_I.branch[9].l_um_iw[202] ;
 wire \top_I.branch[9].l_um_iw[203] ;
 wire \top_I.branch[9].l_um_iw[204] ;
 wire \top_I.branch[9].l_um_iw[205] ;
 wire \top_I.branch[9].l_um_iw[206] ;
 wire \top_I.branch[9].l_um_iw[207] ;
 wire \top_I.branch[9].l_um_iw[208] ;
 wire \top_I.branch[9].l_um_iw[209] ;
 wire \top_I.branch[9].l_um_iw[20] ;
 wire \top_I.branch[9].l_um_iw[210] ;
 wire \top_I.branch[9].l_um_iw[211] ;
 wire \top_I.branch[9].l_um_iw[212] ;
 wire \top_I.branch[9].l_um_iw[213] ;
 wire \top_I.branch[9].l_um_iw[214] ;
 wire \top_I.branch[9].l_um_iw[215] ;
 wire \top_I.branch[9].l_um_iw[216] ;
 wire \top_I.branch[9].l_um_iw[217] ;
 wire \top_I.branch[9].l_um_iw[218] ;
 wire \top_I.branch[9].l_um_iw[219] ;
 wire \top_I.branch[9].l_um_iw[21] ;
 wire \top_I.branch[9].l_um_iw[220] ;
 wire \top_I.branch[9].l_um_iw[221] ;
 wire \top_I.branch[9].l_um_iw[222] ;
 wire \top_I.branch[9].l_um_iw[223] ;
 wire \top_I.branch[9].l_um_iw[224] ;
 wire \top_I.branch[9].l_um_iw[225] ;
 wire \top_I.branch[9].l_um_iw[226] ;
 wire \top_I.branch[9].l_um_iw[227] ;
 wire \top_I.branch[9].l_um_iw[228] ;
 wire \top_I.branch[9].l_um_iw[229] ;
 wire \top_I.branch[9].l_um_iw[22] ;
 wire \top_I.branch[9].l_um_iw[230] ;
 wire \top_I.branch[9].l_um_iw[231] ;
 wire \top_I.branch[9].l_um_iw[232] ;
 wire \top_I.branch[9].l_um_iw[233] ;
 wire \top_I.branch[9].l_um_iw[234] ;
 wire \top_I.branch[9].l_um_iw[235] ;
 wire \top_I.branch[9].l_um_iw[236] ;
 wire \top_I.branch[9].l_um_iw[237] ;
 wire \top_I.branch[9].l_um_iw[238] ;
 wire \top_I.branch[9].l_um_iw[239] ;
 wire \top_I.branch[9].l_um_iw[23] ;
 wire \top_I.branch[9].l_um_iw[240] ;
 wire \top_I.branch[9].l_um_iw[241] ;
 wire \top_I.branch[9].l_um_iw[242] ;
 wire \top_I.branch[9].l_um_iw[243] ;
 wire \top_I.branch[9].l_um_iw[244] ;
 wire \top_I.branch[9].l_um_iw[245] ;
 wire \top_I.branch[9].l_um_iw[246] ;
 wire \top_I.branch[9].l_um_iw[247] ;
 wire \top_I.branch[9].l_um_iw[248] ;
 wire \top_I.branch[9].l_um_iw[249] ;
 wire \top_I.branch[9].l_um_iw[24] ;
 wire \top_I.branch[9].l_um_iw[250] ;
 wire \top_I.branch[9].l_um_iw[251] ;
 wire \top_I.branch[9].l_um_iw[252] ;
 wire \top_I.branch[9].l_um_iw[253] ;
 wire \top_I.branch[9].l_um_iw[254] ;
 wire \top_I.branch[9].l_um_iw[255] ;
 wire \top_I.branch[9].l_um_iw[256] ;
 wire \top_I.branch[9].l_um_iw[257] ;
 wire \top_I.branch[9].l_um_iw[258] ;
 wire \top_I.branch[9].l_um_iw[259] ;
 wire \top_I.branch[9].l_um_iw[25] ;
 wire \top_I.branch[9].l_um_iw[260] ;
 wire \top_I.branch[9].l_um_iw[261] ;
 wire \top_I.branch[9].l_um_iw[262] ;
 wire \top_I.branch[9].l_um_iw[263] ;
 wire \top_I.branch[9].l_um_iw[264] ;
 wire \top_I.branch[9].l_um_iw[265] ;
 wire \top_I.branch[9].l_um_iw[266] ;
 wire \top_I.branch[9].l_um_iw[267] ;
 wire \top_I.branch[9].l_um_iw[268] ;
 wire \top_I.branch[9].l_um_iw[269] ;
 wire \top_I.branch[9].l_um_iw[26] ;
 wire \top_I.branch[9].l_um_iw[270] ;
 wire \top_I.branch[9].l_um_iw[271] ;
 wire \top_I.branch[9].l_um_iw[272] ;
 wire \top_I.branch[9].l_um_iw[273] ;
 wire \top_I.branch[9].l_um_iw[274] ;
 wire \top_I.branch[9].l_um_iw[275] ;
 wire \top_I.branch[9].l_um_iw[276] ;
 wire \top_I.branch[9].l_um_iw[277] ;
 wire \top_I.branch[9].l_um_iw[278] ;
 wire \top_I.branch[9].l_um_iw[279] ;
 wire \top_I.branch[9].l_um_iw[27] ;
 wire \top_I.branch[9].l_um_iw[280] ;
 wire \top_I.branch[9].l_um_iw[281] ;
 wire \top_I.branch[9].l_um_iw[282] ;
 wire \top_I.branch[9].l_um_iw[283] ;
 wire \top_I.branch[9].l_um_iw[284] ;
 wire \top_I.branch[9].l_um_iw[285] ;
 wire \top_I.branch[9].l_um_iw[286] ;
 wire \top_I.branch[9].l_um_iw[287] ;
 wire \top_I.branch[9].l_um_iw[28] ;
 wire \top_I.branch[9].l_um_iw[29] ;
 wire \top_I.branch[9].l_um_iw[2] ;
 wire \top_I.branch[9].l_um_iw[30] ;
 wire \top_I.branch[9].l_um_iw[31] ;
 wire \top_I.branch[9].l_um_iw[32] ;
 wire \top_I.branch[9].l_um_iw[33] ;
 wire \top_I.branch[9].l_um_iw[34] ;
 wire \top_I.branch[9].l_um_iw[35] ;
 wire \top_I.branch[9].l_um_iw[36] ;
 wire \top_I.branch[9].l_um_iw[37] ;
 wire \top_I.branch[9].l_um_iw[38] ;
 wire \top_I.branch[9].l_um_iw[39] ;
 wire \top_I.branch[9].l_um_iw[3] ;
 wire \top_I.branch[9].l_um_iw[40] ;
 wire \top_I.branch[9].l_um_iw[41] ;
 wire \top_I.branch[9].l_um_iw[42] ;
 wire \top_I.branch[9].l_um_iw[43] ;
 wire \top_I.branch[9].l_um_iw[44] ;
 wire \top_I.branch[9].l_um_iw[45] ;
 wire \top_I.branch[9].l_um_iw[46] ;
 wire \top_I.branch[9].l_um_iw[47] ;
 wire \top_I.branch[9].l_um_iw[48] ;
 wire \top_I.branch[9].l_um_iw[49] ;
 wire \top_I.branch[9].l_um_iw[4] ;
 wire \top_I.branch[9].l_um_iw[50] ;
 wire \top_I.branch[9].l_um_iw[51] ;
 wire \top_I.branch[9].l_um_iw[52] ;
 wire \top_I.branch[9].l_um_iw[53] ;
 wire \top_I.branch[9].l_um_iw[54] ;
 wire \top_I.branch[9].l_um_iw[55] ;
 wire \top_I.branch[9].l_um_iw[56] ;
 wire \top_I.branch[9].l_um_iw[57] ;
 wire \top_I.branch[9].l_um_iw[58] ;
 wire \top_I.branch[9].l_um_iw[59] ;
 wire \top_I.branch[9].l_um_iw[5] ;
 wire \top_I.branch[9].l_um_iw[60] ;
 wire \top_I.branch[9].l_um_iw[61] ;
 wire \top_I.branch[9].l_um_iw[62] ;
 wire \top_I.branch[9].l_um_iw[63] ;
 wire \top_I.branch[9].l_um_iw[64] ;
 wire \top_I.branch[9].l_um_iw[65] ;
 wire \top_I.branch[9].l_um_iw[66] ;
 wire \top_I.branch[9].l_um_iw[67] ;
 wire \top_I.branch[9].l_um_iw[68] ;
 wire \top_I.branch[9].l_um_iw[69] ;
 wire \top_I.branch[9].l_um_iw[6] ;
 wire \top_I.branch[9].l_um_iw[70] ;
 wire \top_I.branch[9].l_um_iw[71] ;
 wire \top_I.branch[9].l_um_iw[72] ;
 wire \top_I.branch[9].l_um_iw[73] ;
 wire \top_I.branch[9].l_um_iw[74] ;
 wire \top_I.branch[9].l_um_iw[75] ;
 wire \top_I.branch[9].l_um_iw[76] ;
 wire \top_I.branch[9].l_um_iw[77] ;
 wire \top_I.branch[9].l_um_iw[78] ;
 wire \top_I.branch[9].l_um_iw[79] ;
 wire \top_I.branch[9].l_um_iw[7] ;
 wire \top_I.branch[9].l_um_iw[80] ;
 wire \top_I.branch[9].l_um_iw[81] ;
 wire \top_I.branch[9].l_um_iw[82] ;
 wire \top_I.branch[9].l_um_iw[83] ;
 wire \top_I.branch[9].l_um_iw[84] ;
 wire \top_I.branch[9].l_um_iw[85] ;
 wire \top_I.branch[9].l_um_iw[86] ;
 wire \top_I.branch[9].l_um_iw[87] ;
 wire \top_I.branch[9].l_um_iw[88] ;
 wire \top_I.branch[9].l_um_iw[89] ;
 wire \top_I.branch[9].l_um_iw[8] ;
 wire \top_I.branch[9].l_um_iw[90] ;
 wire \top_I.branch[9].l_um_iw[91] ;
 wire \top_I.branch[9].l_um_iw[92] ;
 wire \top_I.branch[9].l_um_iw[93] ;
 wire \top_I.branch[9].l_um_iw[94] ;
 wire \top_I.branch[9].l_um_iw[95] ;
 wire \top_I.branch[9].l_um_iw[96] ;
 wire \top_I.branch[9].l_um_iw[97] ;
 wire \top_I.branch[9].l_um_iw[98] ;
 wire \top_I.branch[9].l_um_iw[99] ;
 wire \top_I.branch[9].l_um_iw[9] ;
 wire \top_I.branch[9].l_um_k_zero[0] ;
 wire \top_I.branch[9].l_um_k_zero[10] ;
 wire \top_I.branch[9].l_um_k_zero[11] ;
 wire \top_I.branch[9].l_um_k_zero[12] ;
 wire \top_I.branch[9].l_um_k_zero[13] ;
 wire \top_I.branch[9].l_um_k_zero[14] ;
 wire \top_I.branch[9].l_um_k_zero[15] ;
 wire \top_I.branch[9].l_um_k_zero[1] ;
 wire \top_I.branch[9].l_um_k_zero[2] ;
 wire \top_I.branch[9].l_um_k_zero[3] ;
 wire \top_I.branch[9].l_um_k_zero[4] ;
 wire \top_I.branch[9].l_um_k_zero[5] ;
 wire \top_I.branch[9].l_um_k_zero[6] ;
 wire \top_I.branch[9].l_um_k_zero[7] ;
 wire \top_I.branch[9].l_um_k_zero[8] ;
 wire \top_I.branch[9].l_um_k_zero[9] ;
 wire \top_I.k_one ;
 wire \top_I.spine_iw[0] ;
 wire \top_I.spine_iw[10] ;
 wire \top_I.spine_iw[11] ;
 wire \top_I.spine_iw[12] ;
 wire \top_I.spine_iw[13] ;
 wire \top_I.spine_iw[14] ;
 wire \top_I.spine_iw[15] ;
 wire \top_I.spine_iw[16] ;
 wire \top_I.spine_iw[17] ;
 wire \top_I.spine_iw[18] ;
 wire \top_I.spine_iw[19] ;
 wire \top_I.spine_iw[1] ;
 wire \top_I.spine_iw[20] ;
 wire \top_I.spine_iw[21] ;
 wire \top_I.spine_iw[22] ;
 wire \top_I.spine_iw[23] ;
 wire \top_I.spine_iw[24] ;
 wire \top_I.spine_iw[25] ;
 wire \top_I.spine_iw[26] ;
 wire \top_I.spine_iw[27] ;
 wire \top_I.spine_iw[28] ;
 wire \top_I.spine_iw[29] ;
 wire \top_I.spine_iw[2] ;
 wire \top_I.spine_iw[30] ;
 wire \top_I.spine_iw[3] ;
 wire \top_I.spine_iw[4] ;
 wire \top_I.spine_iw[5] ;
 wire \top_I.spine_iw[6] ;
 wire \top_I.spine_iw[7] ;
 wire \top_I.spine_iw[8] ;
 wire \top_I.spine_iw[9] ;
 wire \top_I.spine_ow[0] ;
 wire \top_I.spine_ow[10] ;
 wire \top_I.spine_ow[11] ;
 wire \top_I.spine_ow[12] ;
 wire \top_I.spine_ow[13] ;
 wire \top_I.spine_ow[14] ;
 wire \top_I.spine_ow[15] ;
 wire \top_I.spine_ow[16] ;
 wire \top_I.spine_ow[17] ;
 wire \top_I.spine_ow[18] ;
 wire \top_I.spine_ow[19] ;
 wire \top_I.spine_ow[1] ;
 wire \top_I.spine_ow[20] ;
 wire \top_I.spine_ow[21] ;
 wire \top_I.spine_ow[22] ;
 wire \top_I.spine_ow[23] ;
 wire \top_I.spine_ow[24] ;
 wire \top_I.spine_ow[25] ;
 wire \top_I.spine_ow[2] ;
 wire \top_I.spine_ow[3] ;
 wire \top_I.spine_ow[4] ;
 wire \top_I.spine_ow[5] ;
 wire \top_I.spine_ow[6] ;
 wire \top_I.spine_ow[7] ;
 wire \top_I.spine_ow[8] ;
 wire \top_I.spine_ow[9] ;

 tt_um_loopback \top_I.branch[0].col_um[0].um_bot_I.block_0_0.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[0] ),
    .ena(\top_I.branch[0].l_um_ena[0] ),
    .rst_n(\top_I.branch[0].l_um_iw[1] ),
    .ui_in({\top_I.branch[0].l_um_iw[9] ,
    \top_I.branch[0].l_um_iw[8] ,
    \top_I.branch[0].l_um_iw[7] ,
    \top_I.branch[0].l_um_iw[6] ,
    \top_I.branch[0].l_um_iw[5] ,
    \top_I.branch[0].l_um_iw[4] ,
    \top_I.branch[0].l_um_iw[3] ,
    \top_I.branch[0].l_um_iw[2] }),
    .uio_in({\top_I.branch[0].l_um_iw[17] ,
    \top_I.branch[0].l_um_iw[16] ,
    \top_I.branch[0].l_um_iw[15] ,
    \top_I.branch[0].l_um_iw[14] ,
    \top_I.branch[0].l_um_iw[13] ,
    \top_I.branch[0].l_um_iw[12] ,
    \top_I.branch[0].l_um_iw[11] ,
    \top_I.branch[0].l_um_iw[10] }),
    .uio_oe({\top_I.branch[0].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_as1802 \top_I.branch[0].col_um[0].um_top_I.block_1_0.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[18] ),
    .ena(\top_I.branch[0].l_um_ena[1] ),
    .rst_n(\top_I.branch[0].l_um_iw[19] ),
    .ui_in({\top_I.branch[0].l_um_iw[27] ,
    \top_I.branch[0].l_um_iw[26] ,
    \top_I.branch[0].l_um_iw[25] ,
    \top_I.branch[0].l_um_iw[24] ,
    \top_I.branch[0].l_um_iw[23] ,
    \top_I.branch[0].l_um_iw[22] ,
    \top_I.branch[0].l_um_iw[21] ,
    \top_I.branch[0].l_um_iw[20] }),
    .uio_in({\top_I.branch[0].l_um_iw[35] ,
    \top_I.branch[0].l_um_iw[34] ,
    \top_I.branch[0].l_um_iw[33] ,
    \top_I.branch[0].l_um_iw[32] ,
    \top_I.branch[0].l_um_iw[31] ,
    \top_I.branch[0].l_um_iw[30] ,
    \top_I.branch[0].l_um_iw[29] ,
    \top_I.branch[0].l_um_iw[28] }),
    .uio_oe({\top_I.branch[0].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[0] }));
 tt_um_wokwi_366318576852367361 \top_I.branch[0].col_um[1].um_bot_I.block_0_1.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[36] ),
    .ena(\top_I.branch[0].l_um_ena[2] ),
    .rst_n(\top_I.branch[0].l_um_iw[37] ),
    .ui_in({\top_I.branch[0].l_um_iw[45] ,
    \top_I.branch[0].l_um_iw[44] ,
    \top_I.branch[0].l_um_iw[43] ,
    \top_I.branch[0].l_um_iw[42] ,
    \top_I.branch[0].l_um_iw[41] ,
    \top_I.branch[0].l_um_iw[40] ,
    \top_I.branch[0].l_um_iw[39] ,
    \top_I.branch[0].l_um_iw[38] }),
    .uio_in({\top_I.branch[0].l_um_iw[53] ,
    \top_I.branch[0].l_um_iw[52] ,
    \top_I.branch[0].l_um_iw[51] ,
    \top_I.branch[0].l_um_iw[50] ,
    \top_I.branch[0].l_um_iw[49] ,
    \top_I.branch[0].l_um_iw[48] ,
    \top_I.branch[0].l_um_iw[47] ,
    \top_I.branch[0].l_um_iw[46] }),
    .uio_oe({\top_I.branch[0].col_um[1].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[1].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[1].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[0] }));
 tt_um_moyes0_top_module \top_I.branch[0].col_um[2].um_bot_I.block_0_2.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[72] ),
    .ena(\top_I.branch[0].l_um_ena[4] ),
    .rst_n(\top_I.branch[0].l_um_iw[73] ),
    .ui_in({\top_I.branch[0].l_um_iw[81] ,
    \top_I.branch[0].l_um_iw[80] ,
    \top_I.branch[0].l_um_iw[79] ,
    \top_I.branch[0].l_um_iw[78] ,
    \top_I.branch[0].l_um_iw[77] ,
    \top_I.branch[0].l_um_iw[76] ,
    \top_I.branch[0].l_um_iw[75] ,
    \top_I.branch[0].l_um_iw[74] }),
    .uio_in({\top_I.branch[0].l_um_iw[89] ,
    \top_I.branch[0].l_um_iw[88] ,
    \top_I.branch[0].l_um_iw[87] ,
    \top_I.branch[0].l_um_iw[86] ,
    \top_I.branch[0].l_um_iw[85] ,
    \top_I.branch[0].l_um_iw[84] ,
    \top_I.branch[0].l_um_iw[83] ,
    \top_I.branch[0].l_um_iw[82] }),
    .uio_oe({\top_I.branch[0].col_um[2].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[2].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[2].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[0] }));
 tt_um_TrainLED2_top \top_I.branch[0].col_um[3].um_bot_I.block_0_3.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[108] ),
    .ena(\top_I.branch[0].l_um_ena[6] ),
    .rst_n(\top_I.branch[0].l_um_iw[109] ),
    .ui_in({\top_I.branch[0].l_um_iw[117] ,
    \top_I.branch[0].l_um_iw[116] ,
    \top_I.branch[0].l_um_iw[115] ,
    \top_I.branch[0].l_um_iw[114] ,
    \top_I.branch[0].l_um_iw[113] ,
    \top_I.branch[0].l_um_iw[112] ,
    \top_I.branch[0].l_um_iw[111] ,
    \top_I.branch[0].l_um_iw[110] }),
    .uio_in({\top_I.branch[0].l_um_iw[125] ,
    \top_I.branch[0].l_um_iw[124] ,
    \top_I.branch[0].l_um_iw[123] ,
    \top_I.branch[0].l_um_iw[122] ,
    \top_I.branch[0].l_um_iw[121] ,
    \top_I.branch[0].l_um_iw[120] ,
    \top_I.branch[0].l_um_iw[119] ,
    \top_I.branch[0].l_um_iw[118] }),
    .uio_oe({\top_I.branch[0].col_um[3].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[3].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[3].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[0] }));
 tt_um_ternaryPC_radixconvert \top_I.branch[0].col_um[4].um_bot_I.block_0_4.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[144] ),
    .ena(\top_I.branch[0].l_um_ena[8] ),
    .rst_n(\top_I.branch[0].l_um_iw[145] ),
    .ui_in({\top_I.branch[0].l_um_iw[153] ,
    \top_I.branch[0].l_um_iw[152] ,
    \top_I.branch[0].l_um_iw[151] ,
    \top_I.branch[0].l_um_iw[150] ,
    \top_I.branch[0].l_um_iw[149] ,
    \top_I.branch[0].l_um_iw[148] ,
    \top_I.branch[0].l_um_iw[147] ,
    \top_I.branch[0].l_um_iw[146] }),
    .uio_in({\top_I.branch[0].l_um_iw[161] ,
    \top_I.branch[0].l_um_iw[160] ,
    \top_I.branch[0].l_um_iw[159] ,
    \top_I.branch[0].l_um_iw[158] ,
    \top_I.branch[0].l_um_iw[157] ,
    \top_I.branch[0].l_um_iw[156] ,
    \top_I.branch[0].l_um_iw[155] ,
    \top_I.branch[0].l_um_iw[154] }),
    .uio_oe({\top_I.branch[0].col_um[4].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[4].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[4].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[0] }));
 tt_um_cam \top_I.branch[0].col_um[5].um_bot_I.block_0_5.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[180] ),
    .ena(\top_I.branch[0].l_um_ena[10] ),
    .rst_n(\top_I.branch[0].l_um_iw[181] ),
    .ui_in({\top_I.branch[0].l_um_iw[189] ,
    \top_I.branch[0].l_um_iw[188] ,
    \top_I.branch[0].l_um_iw[187] ,
    \top_I.branch[0].l_um_iw[186] ,
    \top_I.branch[0].l_um_iw[185] ,
    \top_I.branch[0].l_um_iw[184] ,
    \top_I.branch[0].l_um_iw[183] ,
    \top_I.branch[0].l_um_iw[182] }),
    .uio_in({\top_I.branch[0].l_um_iw[197] ,
    \top_I.branch[0].l_um_iw[196] ,
    \top_I.branch[0].l_um_iw[195] ,
    \top_I.branch[0].l_um_iw[194] ,
    \top_I.branch[0].l_um_iw[193] ,
    \top_I.branch[0].l_um_iw[192] ,
    \top_I.branch[0].l_um_iw[191] ,
    \top_I.branch[0].l_um_iw[190] }),
    .uio_oe({\top_I.branch[0].col_um[5].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[5].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[5].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[0] }));
 tt_um_power_test \top_I.branch[0].col_um[6].um_bot_I.block_0_6.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[216] ),
    .ena(\top_I.branch[0].l_um_ena[12] ),
    .rst_n(\top_I.branch[0].l_um_iw[217] ),
    .ui_in({\top_I.branch[0].l_um_iw[225] ,
    \top_I.branch[0].l_um_iw[224] ,
    \top_I.branch[0].l_um_iw[223] ,
    \top_I.branch[0].l_um_iw[222] ,
    \top_I.branch[0].l_um_iw[221] ,
    \top_I.branch[0].l_um_iw[220] ,
    \top_I.branch[0].l_um_iw[219] ,
    \top_I.branch[0].l_um_iw[218] }),
    .uio_in({\top_I.branch[0].l_um_iw[233] ,
    \top_I.branch[0].l_um_iw[232] ,
    \top_I.branch[0].l_um_iw[231] ,
    \top_I.branch[0].l_um_iw[230] ,
    \top_I.branch[0].l_um_iw[229] ,
    \top_I.branch[0].l_um_iw[228] ,
    \top_I.branch[0].l_um_iw[227] ,
    \top_I.branch[0].l_um_iw[226] }),
    .uio_oe({\top_I.branch[0].col_um[6].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[6].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[6].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[0] }));
 tt_um_ringosc_cnt_pfet \top_I.branch[0].col_um[7].um_bot_I.block_0_7.tt_um_I  (.clk(\top_I.branch[0].l_um_iw[252] ),
    .ena(\top_I.branch[0].l_um_ena[14] ),
    .rst_n(\top_I.branch[0].l_um_iw[253] ),
    .ui_in({\top_I.branch[0].l_um_iw[261] ,
    \top_I.branch[0].l_um_iw[260] ,
    \top_I.branch[0].l_um_iw[259] ,
    \top_I.branch[0].l_um_iw[258] ,
    \top_I.branch[0].l_um_iw[257] ,
    \top_I.branch[0].l_um_iw[256] ,
    \top_I.branch[0].l_um_iw[255] ,
    \top_I.branch[0].l_um_iw[254] }),
    .uio_in({\top_I.branch[0].l_um_iw[269] ,
    \top_I.branch[0].l_um_iw[268] ,
    \top_I.branch[0].l_um_iw[267] ,
    \top_I.branch[0].l_um_iw[266] ,
    \top_I.branch[0].l_um_iw[265] ,
    \top_I.branch[0].l_um_iw[264] ,
    \top_I.branch[0].l_um_iw[263] ,
    \top_I.branch[0].l_um_iw[262] }),
    .uio_oe({\top_I.branch[0].col_um[7].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[0].col_um[7].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[0].col_um[7].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[0].mux_I  (.k_one(\top_I.branch[0].l_k_one ),
    .k_zero(\top_I.branch[0].l_k_zero ),
    .addr({\top_I.branch[0].l_k_zero ,
    \top_I.branch[0].l_k_zero ,
    \top_I.branch[0].l_k_zero ,
    \top_I.branch[0].l_k_zero ,
    \top_I.branch[0].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[0].l_um_ena[15] ,
    \top_I.branch[0].l_um_ena[14] ,
    \top_I.branch[0].l_um_ena[13] ,
    \top_I.branch[0].l_um_ena[12] ,
    \top_I.branch[0].l_um_ena[11] ,
    \top_I.branch[0].l_um_ena[10] ,
    \top_I.branch[0].l_um_ena[9] ,
    \top_I.branch[0].l_um_ena[8] ,
    \top_I.branch[0].l_um_ena[7] ,
    \top_I.branch[0].l_um_ena[6] ,
    \top_I.branch[0].l_um_ena[5] ,
    \top_I.branch[0].l_um_ena[4] ,
    \top_I.branch[0].l_um_ena[3] ,
    \top_I.branch[0].l_um_ena[2] ,
    \top_I.branch[0].l_um_ena[1] ,
    \top_I.branch[0].l_um_ena[0] }),
    .um_iw({\top_I.branch[0].l_um_iw[287] ,
    \top_I.branch[0].l_um_iw[286] ,
    \top_I.branch[0].l_um_iw[285] ,
    \top_I.branch[0].l_um_iw[284] ,
    \top_I.branch[0].l_um_iw[283] ,
    \top_I.branch[0].l_um_iw[282] ,
    \top_I.branch[0].l_um_iw[281] ,
    \top_I.branch[0].l_um_iw[280] ,
    \top_I.branch[0].l_um_iw[279] ,
    \top_I.branch[0].l_um_iw[278] ,
    \top_I.branch[0].l_um_iw[277] ,
    \top_I.branch[0].l_um_iw[276] ,
    \top_I.branch[0].l_um_iw[275] ,
    \top_I.branch[0].l_um_iw[274] ,
    \top_I.branch[0].l_um_iw[273] ,
    \top_I.branch[0].l_um_iw[272] ,
    \top_I.branch[0].l_um_iw[271] ,
    \top_I.branch[0].l_um_iw[270] ,
    \top_I.branch[0].l_um_iw[269] ,
    \top_I.branch[0].l_um_iw[268] ,
    \top_I.branch[0].l_um_iw[267] ,
    \top_I.branch[0].l_um_iw[266] ,
    \top_I.branch[0].l_um_iw[265] ,
    \top_I.branch[0].l_um_iw[264] ,
    \top_I.branch[0].l_um_iw[263] ,
    \top_I.branch[0].l_um_iw[262] ,
    \top_I.branch[0].l_um_iw[261] ,
    \top_I.branch[0].l_um_iw[260] ,
    \top_I.branch[0].l_um_iw[259] ,
    \top_I.branch[0].l_um_iw[258] ,
    \top_I.branch[0].l_um_iw[257] ,
    \top_I.branch[0].l_um_iw[256] ,
    \top_I.branch[0].l_um_iw[255] ,
    \top_I.branch[0].l_um_iw[254] ,
    \top_I.branch[0].l_um_iw[253] ,
    \top_I.branch[0].l_um_iw[252] ,
    \top_I.branch[0].l_um_iw[251] ,
    \top_I.branch[0].l_um_iw[250] ,
    \top_I.branch[0].l_um_iw[249] ,
    \top_I.branch[0].l_um_iw[248] ,
    \top_I.branch[0].l_um_iw[247] ,
    \top_I.branch[0].l_um_iw[246] ,
    \top_I.branch[0].l_um_iw[245] ,
    \top_I.branch[0].l_um_iw[244] ,
    \top_I.branch[0].l_um_iw[243] ,
    \top_I.branch[0].l_um_iw[242] ,
    \top_I.branch[0].l_um_iw[241] ,
    \top_I.branch[0].l_um_iw[240] ,
    \top_I.branch[0].l_um_iw[239] ,
    \top_I.branch[0].l_um_iw[238] ,
    \top_I.branch[0].l_um_iw[237] ,
    \top_I.branch[0].l_um_iw[236] ,
    \top_I.branch[0].l_um_iw[235] ,
    \top_I.branch[0].l_um_iw[234] ,
    \top_I.branch[0].l_um_iw[233] ,
    \top_I.branch[0].l_um_iw[232] ,
    \top_I.branch[0].l_um_iw[231] ,
    \top_I.branch[0].l_um_iw[230] ,
    \top_I.branch[0].l_um_iw[229] ,
    \top_I.branch[0].l_um_iw[228] ,
    \top_I.branch[0].l_um_iw[227] ,
    \top_I.branch[0].l_um_iw[226] ,
    \top_I.branch[0].l_um_iw[225] ,
    \top_I.branch[0].l_um_iw[224] ,
    \top_I.branch[0].l_um_iw[223] ,
    \top_I.branch[0].l_um_iw[222] ,
    \top_I.branch[0].l_um_iw[221] ,
    \top_I.branch[0].l_um_iw[220] ,
    \top_I.branch[0].l_um_iw[219] ,
    \top_I.branch[0].l_um_iw[218] ,
    \top_I.branch[0].l_um_iw[217] ,
    \top_I.branch[0].l_um_iw[216] ,
    \top_I.branch[0].l_um_iw[215] ,
    \top_I.branch[0].l_um_iw[214] ,
    \top_I.branch[0].l_um_iw[213] ,
    \top_I.branch[0].l_um_iw[212] ,
    \top_I.branch[0].l_um_iw[211] ,
    \top_I.branch[0].l_um_iw[210] ,
    \top_I.branch[0].l_um_iw[209] ,
    \top_I.branch[0].l_um_iw[208] ,
    \top_I.branch[0].l_um_iw[207] ,
    \top_I.branch[0].l_um_iw[206] ,
    \top_I.branch[0].l_um_iw[205] ,
    \top_I.branch[0].l_um_iw[204] ,
    \top_I.branch[0].l_um_iw[203] ,
    \top_I.branch[0].l_um_iw[202] ,
    \top_I.branch[0].l_um_iw[201] ,
    \top_I.branch[0].l_um_iw[200] ,
    \top_I.branch[0].l_um_iw[199] ,
    \top_I.branch[0].l_um_iw[198] ,
    \top_I.branch[0].l_um_iw[197] ,
    \top_I.branch[0].l_um_iw[196] ,
    \top_I.branch[0].l_um_iw[195] ,
    \top_I.branch[0].l_um_iw[194] ,
    \top_I.branch[0].l_um_iw[193] ,
    \top_I.branch[0].l_um_iw[192] ,
    \top_I.branch[0].l_um_iw[191] ,
    \top_I.branch[0].l_um_iw[190] ,
    \top_I.branch[0].l_um_iw[189] ,
    \top_I.branch[0].l_um_iw[188] ,
    \top_I.branch[0].l_um_iw[187] ,
    \top_I.branch[0].l_um_iw[186] ,
    \top_I.branch[0].l_um_iw[185] ,
    \top_I.branch[0].l_um_iw[184] ,
    \top_I.branch[0].l_um_iw[183] ,
    \top_I.branch[0].l_um_iw[182] ,
    \top_I.branch[0].l_um_iw[181] ,
    \top_I.branch[0].l_um_iw[180] ,
    \top_I.branch[0].l_um_iw[179] ,
    \top_I.branch[0].l_um_iw[178] ,
    \top_I.branch[0].l_um_iw[177] ,
    \top_I.branch[0].l_um_iw[176] ,
    \top_I.branch[0].l_um_iw[175] ,
    \top_I.branch[0].l_um_iw[174] ,
    \top_I.branch[0].l_um_iw[173] ,
    \top_I.branch[0].l_um_iw[172] ,
    \top_I.branch[0].l_um_iw[171] ,
    \top_I.branch[0].l_um_iw[170] ,
    \top_I.branch[0].l_um_iw[169] ,
    \top_I.branch[0].l_um_iw[168] ,
    \top_I.branch[0].l_um_iw[167] ,
    \top_I.branch[0].l_um_iw[166] ,
    \top_I.branch[0].l_um_iw[165] ,
    \top_I.branch[0].l_um_iw[164] ,
    \top_I.branch[0].l_um_iw[163] ,
    \top_I.branch[0].l_um_iw[162] ,
    \top_I.branch[0].l_um_iw[161] ,
    \top_I.branch[0].l_um_iw[160] ,
    \top_I.branch[0].l_um_iw[159] ,
    \top_I.branch[0].l_um_iw[158] ,
    \top_I.branch[0].l_um_iw[157] ,
    \top_I.branch[0].l_um_iw[156] ,
    \top_I.branch[0].l_um_iw[155] ,
    \top_I.branch[0].l_um_iw[154] ,
    \top_I.branch[0].l_um_iw[153] ,
    \top_I.branch[0].l_um_iw[152] ,
    \top_I.branch[0].l_um_iw[151] ,
    \top_I.branch[0].l_um_iw[150] ,
    \top_I.branch[0].l_um_iw[149] ,
    \top_I.branch[0].l_um_iw[148] ,
    \top_I.branch[0].l_um_iw[147] ,
    \top_I.branch[0].l_um_iw[146] ,
    \top_I.branch[0].l_um_iw[145] ,
    \top_I.branch[0].l_um_iw[144] ,
    \top_I.branch[0].l_um_iw[143] ,
    \top_I.branch[0].l_um_iw[142] ,
    \top_I.branch[0].l_um_iw[141] ,
    \top_I.branch[0].l_um_iw[140] ,
    \top_I.branch[0].l_um_iw[139] ,
    \top_I.branch[0].l_um_iw[138] ,
    \top_I.branch[0].l_um_iw[137] ,
    \top_I.branch[0].l_um_iw[136] ,
    \top_I.branch[0].l_um_iw[135] ,
    \top_I.branch[0].l_um_iw[134] ,
    \top_I.branch[0].l_um_iw[133] ,
    \top_I.branch[0].l_um_iw[132] ,
    \top_I.branch[0].l_um_iw[131] ,
    \top_I.branch[0].l_um_iw[130] ,
    \top_I.branch[0].l_um_iw[129] ,
    \top_I.branch[0].l_um_iw[128] ,
    \top_I.branch[0].l_um_iw[127] ,
    \top_I.branch[0].l_um_iw[126] ,
    \top_I.branch[0].l_um_iw[125] ,
    \top_I.branch[0].l_um_iw[124] ,
    \top_I.branch[0].l_um_iw[123] ,
    \top_I.branch[0].l_um_iw[122] ,
    \top_I.branch[0].l_um_iw[121] ,
    \top_I.branch[0].l_um_iw[120] ,
    \top_I.branch[0].l_um_iw[119] ,
    \top_I.branch[0].l_um_iw[118] ,
    \top_I.branch[0].l_um_iw[117] ,
    \top_I.branch[0].l_um_iw[116] ,
    \top_I.branch[0].l_um_iw[115] ,
    \top_I.branch[0].l_um_iw[114] ,
    \top_I.branch[0].l_um_iw[113] ,
    \top_I.branch[0].l_um_iw[112] ,
    \top_I.branch[0].l_um_iw[111] ,
    \top_I.branch[0].l_um_iw[110] ,
    \top_I.branch[0].l_um_iw[109] ,
    \top_I.branch[0].l_um_iw[108] ,
    \top_I.branch[0].l_um_iw[107] ,
    \top_I.branch[0].l_um_iw[106] ,
    \top_I.branch[0].l_um_iw[105] ,
    \top_I.branch[0].l_um_iw[104] ,
    \top_I.branch[0].l_um_iw[103] ,
    \top_I.branch[0].l_um_iw[102] ,
    \top_I.branch[0].l_um_iw[101] ,
    \top_I.branch[0].l_um_iw[100] ,
    \top_I.branch[0].l_um_iw[99] ,
    \top_I.branch[0].l_um_iw[98] ,
    \top_I.branch[0].l_um_iw[97] ,
    \top_I.branch[0].l_um_iw[96] ,
    \top_I.branch[0].l_um_iw[95] ,
    \top_I.branch[0].l_um_iw[94] ,
    \top_I.branch[0].l_um_iw[93] ,
    \top_I.branch[0].l_um_iw[92] ,
    \top_I.branch[0].l_um_iw[91] ,
    \top_I.branch[0].l_um_iw[90] ,
    \top_I.branch[0].l_um_iw[89] ,
    \top_I.branch[0].l_um_iw[88] ,
    \top_I.branch[0].l_um_iw[87] ,
    \top_I.branch[0].l_um_iw[86] ,
    \top_I.branch[0].l_um_iw[85] ,
    \top_I.branch[0].l_um_iw[84] ,
    \top_I.branch[0].l_um_iw[83] ,
    \top_I.branch[0].l_um_iw[82] ,
    \top_I.branch[0].l_um_iw[81] ,
    \top_I.branch[0].l_um_iw[80] ,
    \top_I.branch[0].l_um_iw[79] ,
    \top_I.branch[0].l_um_iw[78] ,
    \top_I.branch[0].l_um_iw[77] ,
    \top_I.branch[0].l_um_iw[76] ,
    \top_I.branch[0].l_um_iw[75] ,
    \top_I.branch[0].l_um_iw[74] ,
    \top_I.branch[0].l_um_iw[73] ,
    \top_I.branch[0].l_um_iw[72] ,
    \top_I.branch[0].l_um_iw[71] ,
    \top_I.branch[0].l_um_iw[70] ,
    \top_I.branch[0].l_um_iw[69] ,
    \top_I.branch[0].l_um_iw[68] ,
    \top_I.branch[0].l_um_iw[67] ,
    \top_I.branch[0].l_um_iw[66] ,
    \top_I.branch[0].l_um_iw[65] ,
    \top_I.branch[0].l_um_iw[64] ,
    \top_I.branch[0].l_um_iw[63] ,
    \top_I.branch[0].l_um_iw[62] ,
    \top_I.branch[0].l_um_iw[61] ,
    \top_I.branch[0].l_um_iw[60] ,
    \top_I.branch[0].l_um_iw[59] ,
    \top_I.branch[0].l_um_iw[58] ,
    \top_I.branch[0].l_um_iw[57] ,
    \top_I.branch[0].l_um_iw[56] ,
    \top_I.branch[0].l_um_iw[55] ,
    \top_I.branch[0].l_um_iw[54] ,
    \top_I.branch[0].l_um_iw[53] ,
    \top_I.branch[0].l_um_iw[52] ,
    \top_I.branch[0].l_um_iw[51] ,
    \top_I.branch[0].l_um_iw[50] ,
    \top_I.branch[0].l_um_iw[49] ,
    \top_I.branch[0].l_um_iw[48] ,
    \top_I.branch[0].l_um_iw[47] ,
    \top_I.branch[0].l_um_iw[46] ,
    \top_I.branch[0].l_um_iw[45] ,
    \top_I.branch[0].l_um_iw[44] ,
    \top_I.branch[0].l_um_iw[43] ,
    \top_I.branch[0].l_um_iw[42] ,
    \top_I.branch[0].l_um_iw[41] ,
    \top_I.branch[0].l_um_iw[40] ,
    \top_I.branch[0].l_um_iw[39] ,
    \top_I.branch[0].l_um_iw[38] ,
    \top_I.branch[0].l_um_iw[37] ,
    \top_I.branch[0].l_um_iw[36] ,
    \top_I.branch[0].l_um_iw[35] ,
    \top_I.branch[0].l_um_iw[34] ,
    \top_I.branch[0].l_um_iw[33] ,
    \top_I.branch[0].l_um_iw[32] ,
    \top_I.branch[0].l_um_iw[31] ,
    \top_I.branch[0].l_um_iw[30] ,
    \top_I.branch[0].l_um_iw[29] ,
    \top_I.branch[0].l_um_iw[28] ,
    \top_I.branch[0].l_um_iw[27] ,
    \top_I.branch[0].l_um_iw[26] ,
    \top_I.branch[0].l_um_iw[25] ,
    \top_I.branch[0].l_um_iw[24] ,
    \top_I.branch[0].l_um_iw[23] ,
    \top_I.branch[0].l_um_iw[22] ,
    \top_I.branch[0].l_um_iw[21] ,
    \top_I.branch[0].l_um_iw[20] ,
    \top_I.branch[0].l_um_iw[19] ,
    \top_I.branch[0].l_um_iw[18] ,
    \top_I.branch[0].l_um_iw[17] ,
    \top_I.branch[0].l_um_iw[16] ,
    \top_I.branch[0].l_um_iw[15] ,
    \top_I.branch[0].l_um_iw[14] ,
    \top_I.branch[0].l_um_iw[13] ,
    \top_I.branch[0].l_um_iw[12] ,
    \top_I.branch[0].l_um_iw[11] ,
    \top_I.branch[0].l_um_iw[10] ,
    \top_I.branch[0].l_um_iw[9] ,
    \top_I.branch[0].l_um_iw[8] ,
    \top_I.branch[0].l_um_iw[7] ,
    \top_I.branch[0].l_um_iw[6] ,
    \top_I.branch[0].l_um_iw[5] ,
    \top_I.branch[0].l_um_iw[4] ,
    \top_I.branch[0].l_um_iw[3] ,
    \top_I.branch[0].l_um_iw[2] ,
    \top_I.branch[0].l_um_iw[1] ,
    \top_I.branch[0].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[14] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[12] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[10] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[8] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[6] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[4] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[2] ,
    \top_I.branch[0].l_um_k_zero[1] ,
    \top_I.branch[0].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].l_um_k_zero[15] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[7].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].l_um_k_zero[13] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[6].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].l_um_k_zero[11] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[5].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].l_um_k_zero[9] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[4].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].l_um_k_zero[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[3].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].l_um_k_zero[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[2].um_bot_I.uo_out[0] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].l_um_k_zero[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[1].um_bot_I.uo_out[0] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[0].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[0].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[10].col_um[0].um_top_I.block_11_0.tt_um_I  (.clk(\top_I.branch[10].l_um_iw[18] ),
    .ena(\top_I.branch[10].l_um_ena[1] ),
    .rst_n(\top_I.branch[10].l_um_iw[19] ),
    .ui_in({\top_I.branch[10].l_um_iw[27] ,
    \top_I.branch[10].l_um_iw[26] ,
    \top_I.branch[10].l_um_iw[25] ,
    \top_I.branch[10].l_um_iw[24] ,
    \top_I.branch[10].l_um_iw[23] ,
    \top_I.branch[10].l_um_iw[22] ,
    \top_I.branch[10].l_um_iw[21] ,
    \top_I.branch[10].l_um_iw[20] }),
    .uio_in({\top_I.branch[10].l_um_iw[35] ,
    \top_I.branch[10].l_um_iw[34] ,
    \top_I.branch[10].l_um_iw[33] ,
    \top_I.branch[10].l_um_iw[32] ,
    \top_I.branch[10].l_um_iw[31] ,
    \top_I.branch[10].l_um_iw[30] ,
    \top_I.branch[10].l_um_iw[29] ,
    \top_I.branch[10].l_um_iw[28] }),
    .uio_oe({\top_I.branch[10].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[10].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[10].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[10].mux_I  (.k_one(\top_I.branch[10].l_k_one ),
    .k_zero(\top_I.branch[10].l_k_zero ),
    .addr({\top_I.branch[10].l_k_zero ,
    \top_I.branch[10].l_k_one ,
    \top_I.branch[10].l_k_zero ,
    \top_I.branch[10].l_k_one ,
    \top_I.branch[10].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[10].l_um_ena[15] ,
    \top_I.branch[10].l_um_ena[14] ,
    \top_I.branch[10].l_um_ena[13] ,
    \top_I.branch[10].l_um_ena[12] ,
    \top_I.branch[10].l_um_ena[11] ,
    \top_I.branch[10].l_um_ena[10] ,
    \top_I.branch[10].l_um_ena[9] ,
    \top_I.branch[10].l_um_ena[8] ,
    \top_I.branch[10].l_um_ena[7] ,
    \top_I.branch[10].l_um_ena[6] ,
    \top_I.branch[10].l_um_ena[5] ,
    \top_I.branch[10].l_um_ena[4] ,
    \top_I.branch[10].l_um_ena[3] ,
    \top_I.branch[10].l_um_ena[2] ,
    \top_I.branch[10].l_um_ena[1] ,
    \top_I.branch[10].l_um_ena[0] }),
    .um_iw({\top_I.branch[10].l_um_iw[287] ,
    \top_I.branch[10].l_um_iw[286] ,
    \top_I.branch[10].l_um_iw[285] ,
    \top_I.branch[10].l_um_iw[284] ,
    \top_I.branch[10].l_um_iw[283] ,
    \top_I.branch[10].l_um_iw[282] ,
    \top_I.branch[10].l_um_iw[281] ,
    \top_I.branch[10].l_um_iw[280] ,
    \top_I.branch[10].l_um_iw[279] ,
    \top_I.branch[10].l_um_iw[278] ,
    \top_I.branch[10].l_um_iw[277] ,
    \top_I.branch[10].l_um_iw[276] ,
    \top_I.branch[10].l_um_iw[275] ,
    \top_I.branch[10].l_um_iw[274] ,
    \top_I.branch[10].l_um_iw[273] ,
    \top_I.branch[10].l_um_iw[272] ,
    \top_I.branch[10].l_um_iw[271] ,
    \top_I.branch[10].l_um_iw[270] ,
    \top_I.branch[10].l_um_iw[269] ,
    \top_I.branch[10].l_um_iw[268] ,
    \top_I.branch[10].l_um_iw[267] ,
    \top_I.branch[10].l_um_iw[266] ,
    \top_I.branch[10].l_um_iw[265] ,
    \top_I.branch[10].l_um_iw[264] ,
    \top_I.branch[10].l_um_iw[263] ,
    \top_I.branch[10].l_um_iw[262] ,
    \top_I.branch[10].l_um_iw[261] ,
    \top_I.branch[10].l_um_iw[260] ,
    \top_I.branch[10].l_um_iw[259] ,
    \top_I.branch[10].l_um_iw[258] ,
    \top_I.branch[10].l_um_iw[257] ,
    \top_I.branch[10].l_um_iw[256] ,
    \top_I.branch[10].l_um_iw[255] ,
    \top_I.branch[10].l_um_iw[254] ,
    \top_I.branch[10].l_um_iw[253] ,
    \top_I.branch[10].l_um_iw[252] ,
    \top_I.branch[10].l_um_iw[251] ,
    \top_I.branch[10].l_um_iw[250] ,
    \top_I.branch[10].l_um_iw[249] ,
    \top_I.branch[10].l_um_iw[248] ,
    \top_I.branch[10].l_um_iw[247] ,
    \top_I.branch[10].l_um_iw[246] ,
    \top_I.branch[10].l_um_iw[245] ,
    \top_I.branch[10].l_um_iw[244] ,
    \top_I.branch[10].l_um_iw[243] ,
    \top_I.branch[10].l_um_iw[242] ,
    \top_I.branch[10].l_um_iw[241] ,
    \top_I.branch[10].l_um_iw[240] ,
    \top_I.branch[10].l_um_iw[239] ,
    \top_I.branch[10].l_um_iw[238] ,
    \top_I.branch[10].l_um_iw[237] ,
    \top_I.branch[10].l_um_iw[236] ,
    \top_I.branch[10].l_um_iw[235] ,
    \top_I.branch[10].l_um_iw[234] ,
    \top_I.branch[10].l_um_iw[233] ,
    \top_I.branch[10].l_um_iw[232] ,
    \top_I.branch[10].l_um_iw[231] ,
    \top_I.branch[10].l_um_iw[230] ,
    \top_I.branch[10].l_um_iw[229] ,
    \top_I.branch[10].l_um_iw[228] ,
    \top_I.branch[10].l_um_iw[227] ,
    \top_I.branch[10].l_um_iw[226] ,
    \top_I.branch[10].l_um_iw[225] ,
    \top_I.branch[10].l_um_iw[224] ,
    \top_I.branch[10].l_um_iw[223] ,
    \top_I.branch[10].l_um_iw[222] ,
    \top_I.branch[10].l_um_iw[221] ,
    \top_I.branch[10].l_um_iw[220] ,
    \top_I.branch[10].l_um_iw[219] ,
    \top_I.branch[10].l_um_iw[218] ,
    \top_I.branch[10].l_um_iw[217] ,
    \top_I.branch[10].l_um_iw[216] ,
    \top_I.branch[10].l_um_iw[215] ,
    \top_I.branch[10].l_um_iw[214] ,
    \top_I.branch[10].l_um_iw[213] ,
    \top_I.branch[10].l_um_iw[212] ,
    \top_I.branch[10].l_um_iw[211] ,
    \top_I.branch[10].l_um_iw[210] ,
    \top_I.branch[10].l_um_iw[209] ,
    \top_I.branch[10].l_um_iw[208] ,
    \top_I.branch[10].l_um_iw[207] ,
    \top_I.branch[10].l_um_iw[206] ,
    \top_I.branch[10].l_um_iw[205] ,
    \top_I.branch[10].l_um_iw[204] ,
    \top_I.branch[10].l_um_iw[203] ,
    \top_I.branch[10].l_um_iw[202] ,
    \top_I.branch[10].l_um_iw[201] ,
    \top_I.branch[10].l_um_iw[200] ,
    \top_I.branch[10].l_um_iw[199] ,
    \top_I.branch[10].l_um_iw[198] ,
    \top_I.branch[10].l_um_iw[197] ,
    \top_I.branch[10].l_um_iw[196] ,
    \top_I.branch[10].l_um_iw[195] ,
    \top_I.branch[10].l_um_iw[194] ,
    \top_I.branch[10].l_um_iw[193] ,
    \top_I.branch[10].l_um_iw[192] ,
    \top_I.branch[10].l_um_iw[191] ,
    \top_I.branch[10].l_um_iw[190] ,
    \top_I.branch[10].l_um_iw[189] ,
    \top_I.branch[10].l_um_iw[188] ,
    \top_I.branch[10].l_um_iw[187] ,
    \top_I.branch[10].l_um_iw[186] ,
    \top_I.branch[10].l_um_iw[185] ,
    \top_I.branch[10].l_um_iw[184] ,
    \top_I.branch[10].l_um_iw[183] ,
    \top_I.branch[10].l_um_iw[182] ,
    \top_I.branch[10].l_um_iw[181] ,
    \top_I.branch[10].l_um_iw[180] ,
    \top_I.branch[10].l_um_iw[179] ,
    \top_I.branch[10].l_um_iw[178] ,
    \top_I.branch[10].l_um_iw[177] ,
    \top_I.branch[10].l_um_iw[176] ,
    \top_I.branch[10].l_um_iw[175] ,
    \top_I.branch[10].l_um_iw[174] ,
    \top_I.branch[10].l_um_iw[173] ,
    \top_I.branch[10].l_um_iw[172] ,
    \top_I.branch[10].l_um_iw[171] ,
    \top_I.branch[10].l_um_iw[170] ,
    \top_I.branch[10].l_um_iw[169] ,
    \top_I.branch[10].l_um_iw[168] ,
    \top_I.branch[10].l_um_iw[167] ,
    \top_I.branch[10].l_um_iw[166] ,
    \top_I.branch[10].l_um_iw[165] ,
    \top_I.branch[10].l_um_iw[164] ,
    \top_I.branch[10].l_um_iw[163] ,
    \top_I.branch[10].l_um_iw[162] ,
    \top_I.branch[10].l_um_iw[161] ,
    \top_I.branch[10].l_um_iw[160] ,
    \top_I.branch[10].l_um_iw[159] ,
    \top_I.branch[10].l_um_iw[158] ,
    \top_I.branch[10].l_um_iw[157] ,
    \top_I.branch[10].l_um_iw[156] ,
    \top_I.branch[10].l_um_iw[155] ,
    \top_I.branch[10].l_um_iw[154] ,
    \top_I.branch[10].l_um_iw[153] ,
    \top_I.branch[10].l_um_iw[152] ,
    \top_I.branch[10].l_um_iw[151] ,
    \top_I.branch[10].l_um_iw[150] ,
    \top_I.branch[10].l_um_iw[149] ,
    \top_I.branch[10].l_um_iw[148] ,
    \top_I.branch[10].l_um_iw[147] ,
    \top_I.branch[10].l_um_iw[146] ,
    \top_I.branch[10].l_um_iw[145] ,
    \top_I.branch[10].l_um_iw[144] ,
    \top_I.branch[10].l_um_iw[143] ,
    \top_I.branch[10].l_um_iw[142] ,
    \top_I.branch[10].l_um_iw[141] ,
    \top_I.branch[10].l_um_iw[140] ,
    \top_I.branch[10].l_um_iw[139] ,
    \top_I.branch[10].l_um_iw[138] ,
    \top_I.branch[10].l_um_iw[137] ,
    \top_I.branch[10].l_um_iw[136] ,
    \top_I.branch[10].l_um_iw[135] ,
    \top_I.branch[10].l_um_iw[134] ,
    \top_I.branch[10].l_um_iw[133] ,
    \top_I.branch[10].l_um_iw[132] ,
    \top_I.branch[10].l_um_iw[131] ,
    \top_I.branch[10].l_um_iw[130] ,
    \top_I.branch[10].l_um_iw[129] ,
    \top_I.branch[10].l_um_iw[128] ,
    \top_I.branch[10].l_um_iw[127] ,
    \top_I.branch[10].l_um_iw[126] ,
    \top_I.branch[10].l_um_iw[125] ,
    \top_I.branch[10].l_um_iw[124] ,
    \top_I.branch[10].l_um_iw[123] ,
    \top_I.branch[10].l_um_iw[122] ,
    \top_I.branch[10].l_um_iw[121] ,
    \top_I.branch[10].l_um_iw[120] ,
    \top_I.branch[10].l_um_iw[119] ,
    \top_I.branch[10].l_um_iw[118] ,
    \top_I.branch[10].l_um_iw[117] ,
    \top_I.branch[10].l_um_iw[116] ,
    \top_I.branch[10].l_um_iw[115] ,
    \top_I.branch[10].l_um_iw[114] ,
    \top_I.branch[10].l_um_iw[113] ,
    \top_I.branch[10].l_um_iw[112] ,
    \top_I.branch[10].l_um_iw[111] ,
    \top_I.branch[10].l_um_iw[110] ,
    \top_I.branch[10].l_um_iw[109] ,
    \top_I.branch[10].l_um_iw[108] ,
    \top_I.branch[10].l_um_iw[107] ,
    \top_I.branch[10].l_um_iw[106] ,
    \top_I.branch[10].l_um_iw[105] ,
    \top_I.branch[10].l_um_iw[104] ,
    \top_I.branch[10].l_um_iw[103] ,
    \top_I.branch[10].l_um_iw[102] ,
    \top_I.branch[10].l_um_iw[101] ,
    \top_I.branch[10].l_um_iw[100] ,
    \top_I.branch[10].l_um_iw[99] ,
    \top_I.branch[10].l_um_iw[98] ,
    \top_I.branch[10].l_um_iw[97] ,
    \top_I.branch[10].l_um_iw[96] ,
    \top_I.branch[10].l_um_iw[95] ,
    \top_I.branch[10].l_um_iw[94] ,
    \top_I.branch[10].l_um_iw[93] ,
    \top_I.branch[10].l_um_iw[92] ,
    \top_I.branch[10].l_um_iw[91] ,
    \top_I.branch[10].l_um_iw[90] ,
    \top_I.branch[10].l_um_iw[89] ,
    \top_I.branch[10].l_um_iw[88] ,
    \top_I.branch[10].l_um_iw[87] ,
    \top_I.branch[10].l_um_iw[86] ,
    \top_I.branch[10].l_um_iw[85] ,
    \top_I.branch[10].l_um_iw[84] ,
    \top_I.branch[10].l_um_iw[83] ,
    \top_I.branch[10].l_um_iw[82] ,
    \top_I.branch[10].l_um_iw[81] ,
    \top_I.branch[10].l_um_iw[80] ,
    \top_I.branch[10].l_um_iw[79] ,
    \top_I.branch[10].l_um_iw[78] ,
    \top_I.branch[10].l_um_iw[77] ,
    \top_I.branch[10].l_um_iw[76] ,
    \top_I.branch[10].l_um_iw[75] ,
    \top_I.branch[10].l_um_iw[74] ,
    \top_I.branch[10].l_um_iw[73] ,
    \top_I.branch[10].l_um_iw[72] ,
    \top_I.branch[10].l_um_iw[71] ,
    \top_I.branch[10].l_um_iw[70] ,
    \top_I.branch[10].l_um_iw[69] ,
    \top_I.branch[10].l_um_iw[68] ,
    \top_I.branch[10].l_um_iw[67] ,
    \top_I.branch[10].l_um_iw[66] ,
    \top_I.branch[10].l_um_iw[65] ,
    \top_I.branch[10].l_um_iw[64] ,
    \top_I.branch[10].l_um_iw[63] ,
    \top_I.branch[10].l_um_iw[62] ,
    \top_I.branch[10].l_um_iw[61] ,
    \top_I.branch[10].l_um_iw[60] ,
    \top_I.branch[10].l_um_iw[59] ,
    \top_I.branch[10].l_um_iw[58] ,
    \top_I.branch[10].l_um_iw[57] ,
    \top_I.branch[10].l_um_iw[56] ,
    \top_I.branch[10].l_um_iw[55] ,
    \top_I.branch[10].l_um_iw[54] ,
    \top_I.branch[10].l_um_iw[53] ,
    \top_I.branch[10].l_um_iw[52] ,
    \top_I.branch[10].l_um_iw[51] ,
    \top_I.branch[10].l_um_iw[50] ,
    \top_I.branch[10].l_um_iw[49] ,
    \top_I.branch[10].l_um_iw[48] ,
    \top_I.branch[10].l_um_iw[47] ,
    \top_I.branch[10].l_um_iw[46] ,
    \top_I.branch[10].l_um_iw[45] ,
    \top_I.branch[10].l_um_iw[44] ,
    \top_I.branch[10].l_um_iw[43] ,
    \top_I.branch[10].l_um_iw[42] ,
    \top_I.branch[10].l_um_iw[41] ,
    \top_I.branch[10].l_um_iw[40] ,
    \top_I.branch[10].l_um_iw[39] ,
    \top_I.branch[10].l_um_iw[38] ,
    \top_I.branch[10].l_um_iw[37] ,
    \top_I.branch[10].l_um_iw[36] ,
    \top_I.branch[10].l_um_iw[35] ,
    \top_I.branch[10].l_um_iw[34] ,
    \top_I.branch[10].l_um_iw[33] ,
    \top_I.branch[10].l_um_iw[32] ,
    \top_I.branch[10].l_um_iw[31] ,
    \top_I.branch[10].l_um_iw[30] ,
    \top_I.branch[10].l_um_iw[29] ,
    \top_I.branch[10].l_um_iw[28] ,
    \top_I.branch[10].l_um_iw[27] ,
    \top_I.branch[10].l_um_iw[26] ,
    \top_I.branch[10].l_um_iw[25] ,
    \top_I.branch[10].l_um_iw[24] ,
    \top_I.branch[10].l_um_iw[23] ,
    \top_I.branch[10].l_um_iw[22] ,
    \top_I.branch[10].l_um_iw[21] ,
    \top_I.branch[10].l_um_iw[20] ,
    \top_I.branch[10].l_um_iw[19] ,
    \top_I.branch[10].l_um_iw[18] ,
    \top_I.branch[10].l_um_iw[17] ,
    \top_I.branch[10].l_um_iw[16] ,
    \top_I.branch[10].l_um_iw[15] ,
    \top_I.branch[10].l_um_iw[14] ,
    \top_I.branch[10].l_um_iw[13] ,
    \top_I.branch[10].l_um_iw[12] ,
    \top_I.branch[10].l_um_iw[11] ,
    \top_I.branch[10].l_um_iw[10] ,
    \top_I.branch[10].l_um_iw[9] ,
    \top_I.branch[10].l_um_iw[8] ,
    \top_I.branch[10].l_um_iw[7] ,
    \top_I.branch[10].l_um_iw[6] ,
    \top_I.branch[10].l_um_iw[5] ,
    \top_I.branch[10].l_um_iw[4] ,
    \top_I.branch[10].l_um_iw[3] ,
    \top_I.branch[10].l_um_iw[2] ,
    \top_I.branch[10].l_um_iw[1] ,
    \top_I.branch[10].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[1] ,
    \top_I.branch[10].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[15] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[14] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[13] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[12] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[11] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[10] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[9] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[8] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[7] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[6] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[5] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[4] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[3] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].l_um_k_zero[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[10].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] ,
    \top_I.branch[10].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[11].col_um[0].um_top_I.block_11_16.tt_um_I  (.clk(\top_I.branch[11].l_um_iw[18] ),
    .ena(\top_I.branch[11].l_um_ena[1] ),
    .rst_n(\top_I.branch[11].l_um_iw[19] ),
    .ui_in({\top_I.branch[11].l_um_iw[27] ,
    \top_I.branch[11].l_um_iw[26] ,
    \top_I.branch[11].l_um_iw[25] ,
    \top_I.branch[11].l_um_iw[24] ,
    \top_I.branch[11].l_um_iw[23] ,
    \top_I.branch[11].l_um_iw[22] ,
    \top_I.branch[11].l_um_iw[21] ,
    \top_I.branch[11].l_um_iw[20] }),
    .uio_in({\top_I.branch[11].l_um_iw[35] ,
    \top_I.branch[11].l_um_iw[34] ,
    \top_I.branch[11].l_um_iw[33] ,
    \top_I.branch[11].l_um_iw[32] ,
    \top_I.branch[11].l_um_iw[31] ,
    \top_I.branch[11].l_um_iw[30] ,
    \top_I.branch[11].l_um_iw[29] ,
    \top_I.branch[11].l_um_iw[28] }),
    .uio_oe({\top_I.branch[11].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[11].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[11].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[11].mux_I  (.k_one(\top_I.branch[11].l_k_one ),
    .k_zero(\top_I.branch[11].l_k_zero ),
    .addr({\top_I.branch[11].l_k_zero ,
    \top_I.branch[11].l_k_one ,
    \top_I.branch[11].l_k_zero ,
    \top_I.branch[11].l_k_one ,
    \top_I.branch[11].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[11].l_um_ena[15] ,
    \top_I.branch[11].l_um_ena[14] ,
    \top_I.branch[11].l_um_ena[13] ,
    \top_I.branch[11].l_um_ena[12] ,
    \top_I.branch[11].l_um_ena[11] ,
    \top_I.branch[11].l_um_ena[10] ,
    \top_I.branch[11].l_um_ena[9] ,
    \top_I.branch[11].l_um_ena[8] ,
    \top_I.branch[11].l_um_ena[7] ,
    \top_I.branch[11].l_um_ena[6] ,
    \top_I.branch[11].l_um_ena[5] ,
    \top_I.branch[11].l_um_ena[4] ,
    \top_I.branch[11].l_um_ena[3] ,
    \top_I.branch[11].l_um_ena[2] ,
    \top_I.branch[11].l_um_ena[1] ,
    \top_I.branch[11].l_um_ena[0] }),
    .um_iw({\top_I.branch[11].l_um_iw[287] ,
    \top_I.branch[11].l_um_iw[286] ,
    \top_I.branch[11].l_um_iw[285] ,
    \top_I.branch[11].l_um_iw[284] ,
    \top_I.branch[11].l_um_iw[283] ,
    \top_I.branch[11].l_um_iw[282] ,
    \top_I.branch[11].l_um_iw[281] ,
    \top_I.branch[11].l_um_iw[280] ,
    \top_I.branch[11].l_um_iw[279] ,
    \top_I.branch[11].l_um_iw[278] ,
    \top_I.branch[11].l_um_iw[277] ,
    \top_I.branch[11].l_um_iw[276] ,
    \top_I.branch[11].l_um_iw[275] ,
    \top_I.branch[11].l_um_iw[274] ,
    \top_I.branch[11].l_um_iw[273] ,
    \top_I.branch[11].l_um_iw[272] ,
    \top_I.branch[11].l_um_iw[271] ,
    \top_I.branch[11].l_um_iw[270] ,
    \top_I.branch[11].l_um_iw[269] ,
    \top_I.branch[11].l_um_iw[268] ,
    \top_I.branch[11].l_um_iw[267] ,
    \top_I.branch[11].l_um_iw[266] ,
    \top_I.branch[11].l_um_iw[265] ,
    \top_I.branch[11].l_um_iw[264] ,
    \top_I.branch[11].l_um_iw[263] ,
    \top_I.branch[11].l_um_iw[262] ,
    \top_I.branch[11].l_um_iw[261] ,
    \top_I.branch[11].l_um_iw[260] ,
    \top_I.branch[11].l_um_iw[259] ,
    \top_I.branch[11].l_um_iw[258] ,
    \top_I.branch[11].l_um_iw[257] ,
    \top_I.branch[11].l_um_iw[256] ,
    \top_I.branch[11].l_um_iw[255] ,
    \top_I.branch[11].l_um_iw[254] ,
    \top_I.branch[11].l_um_iw[253] ,
    \top_I.branch[11].l_um_iw[252] ,
    \top_I.branch[11].l_um_iw[251] ,
    \top_I.branch[11].l_um_iw[250] ,
    \top_I.branch[11].l_um_iw[249] ,
    \top_I.branch[11].l_um_iw[248] ,
    \top_I.branch[11].l_um_iw[247] ,
    \top_I.branch[11].l_um_iw[246] ,
    \top_I.branch[11].l_um_iw[245] ,
    \top_I.branch[11].l_um_iw[244] ,
    \top_I.branch[11].l_um_iw[243] ,
    \top_I.branch[11].l_um_iw[242] ,
    \top_I.branch[11].l_um_iw[241] ,
    \top_I.branch[11].l_um_iw[240] ,
    \top_I.branch[11].l_um_iw[239] ,
    \top_I.branch[11].l_um_iw[238] ,
    \top_I.branch[11].l_um_iw[237] ,
    \top_I.branch[11].l_um_iw[236] ,
    \top_I.branch[11].l_um_iw[235] ,
    \top_I.branch[11].l_um_iw[234] ,
    \top_I.branch[11].l_um_iw[233] ,
    \top_I.branch[11].l_um_iw[232] ,
    \top_I.branch[11].l_um_iw[231] ,
    \top_I.branch[11].l_um_iw[230] ,
    \top_I.branch[11].l_um_iw[229] ,
    \top_I.branch[11].l_um_iw[228] ,
    \top_I.branch[11].l_um_iw[227] ,
    \top_I.branch[11].l_um_iw[226] ,
    \top_I.branch[11].l_um_iw[225] ,
    \top_I.branch[11].l_um_iw[224] ,
    \top_I.branch[11].l_um_iw[223] ,
    \top_I.branch[11].l_um_iw[222] ,
    \top_I.branch[11].l_um_iw[221] ,
    \top_I.branch[11].l_um_iw[220] ,
    \top_I.branch[11].l_um_iw[219] ,
    \top_I.branch[11].l_um_iw[218] ,
    \top_I.branch[11].l_um_iw[217] ,
    \top_I.branch[11].l_um_iw[216] ,
    \top_I.branch[11].l_um_iw[215] ,
    \top_I.branch[11].l_um_iw[214] ,
    \top_I.branch[11].l_um_iw[213] ,
    \top_I.branch[11].l_um_iw[212] ,
    \top_I.branch[11].l_um_iw[211] ,
    \top_I.branch[11].l_um_iw[210] ,
    \top_I.branch[11].l_um_iw[209] ,
    \top_I.branch[11].l_um_iw[208] ,
    \top_I.branch[11].l_um_iw[207] ,
    \top_I.branch[11].l_um_iw[206] ,
    \top_I.branch[11].l_um_iw[205] ,
    \top_I.branch[11].l_um_iw[204] ,
    \top_I.branch[11].l_um_iw[203] ,
    \top_I.branch[11].l_um_iw[202] ,
    \top_I.branch[11].l_um_iw[201] ,
    \top_I.branch[11].l_um_iw[200] ,
    \top_I.branch[11].l_um_iw[199] ,
    \top_I.branch[11].l_um_iw[198] ,
    \top_I.branch[11].l_um_iw[197] ,
    \top_I.branch[11].l_um_iw[196] ,
    \top_I.branch[11].l_um_iw[195] ,
    \top_I.branch[11].l_um_iw[194] ,
    \top_I.branch[11].l_um_iw[193] ,
    \top_I.branch[11].l_um_iw[192] ,
    \top_I.branch[11].l_um_iw[191] ,
    \top_I.branch[11].l_um_iw[190] ,
    \top_I.branch[11].l_um_iw[189] ,
    \top_I.branch[11].l_um_iw[188] ,
    \top_I.branch[11].l_um_iw[187] ,
    \top_I.branch[11].l_um_iw[186] ,
    \top_I.branch[11].l_um_iw[185] ,
    \top_I.branch[11].l_um_iw[184] ,
    \top_I.branch[11].l_um_iw[183] ,
    \top_I.branch[11].l_um_iw[182] ,
    \top_I.branch[11].l_um_iw[181] ,
    \top_I.branch[11].l_um_iw[180] ,
    \top_I.branch[11].l_um_iw[179] ,
    \top_I.branch[11].l_um_iw[178] ,
    \top_I.branch[11].l_um_iw[177] ,
    \top_I.branch[11].l_um_iw[176] ,
    \top_I.branch[11].l_um_iw[175] ,
    \top_I.branch[11].l_um_iw[174] ,
    \top_I.branch[11].l_um_iw[173] ,
    \top_I.branch[11].l_um_iw[172] ,
    \top_I.branch[11].l_um_iw[171] ,
    \top_I.branch[11].l_um_iw[170] ,
    \top_I.branch[11].l_um_iw[169] ,
    \top_I.branch[11].l_um_iw[168] ,
    \top_I.branch[11].l_um_iw[167] ,
    \top_I.branch[11].l_um_iw[166] ,
    \top_I.branch[11].l_um_iw[165] ,
    \top_I.branch[11].l_um_iw[164] ,
    \top_I.branch[11].l_um_iw[163] ,
    \top_I.branch[11].l_um_iw[162] ,
    \top_I.branch[11].l_um_iw[161] ,
    \top_I.branch[11].l_um_iw[160] ,
    \top_I.branch[11].l_um_iw[159] ,
    \top_I.branch[11].l_um_iw[158] ,
    \top_I.branch[11].l_um_iw[157] ,
    \top_I.branch[11].l_um_iw[156] ,
    \top_I.branch[11].l_um_iw[155] ,
    \top_I.branch[11].l_um_iw[154] ,
    \top_I.branch[11].l_um_iw[153] ,
    \top_I.branch[11].l_um_iw[152] ,
    \top_I.branch[11].l_um_iw[151] ,
    \top_I.branch[11].l_um_iw[150] ,
    \top_I.branch[11].l_um_iw[149] ,
    \top_I.branch[11].l_um_iw[148] ,
    \top_I.branch[11].l_um_iw[147] ,
    \top_I.branch[11].l_um_iw[146] ,
    \top_I.branch[11].l_um_iw[145] ,
    \top_I.branch[11].l_um_iw[144] ,
    \top_I.branch[11].l_um_iw[143] ,
    \top_I.branch[11].l_um_iw[142] ,
    \top_I.branch[11].l_um_iw[141] ,
    \top_I.branch[11].l_um_iw[140] ,
    \top_I.branch[11].l_um_iw[139] ,
    \top_I.branch[11].l_um_iw[138] ,
    \top_I.branch[11].l_um_iw[137] ,
    \top_I.branch[11].l_um_iw[136] ,
    \top_I.branch[11].l_um_iw[135] ,
    \top_I.branch[11].l_um_iw[134] ,
    \top_I.branch[11].l_um_iw[133] ,
    \top_I.branch[11].l_um_iw[132] ,
    \top_I.branch[11].l_um_iw[131] ,
    \top_I.branch[11].l_um_iw[130] ,
    \top_I.branch[11].l_um_iw[129] ,
    \top_I.branch[11].l_um_iw[128] ,
    \top_I.branch[11].l_um_iw[127] ,
    \top_I.branch[11].l_um_iw[126] ,
    \top_I.branch[11].l_um_iw[125] ,
    \top_I.branch[11].l_um_iw[124] ,
    \top_I.branch[11].l_um_iw[123] ,
    \top_I.branch[11].l_um_iw[122] ,
    \top_I.branch[11].l_um_iw[121] ,
    \top_I.branch[11].l_um_iw[120] ,
    \top_I.branch[11].l_um_iw[119] ,
    \top_I.branch[11].l_um_iw[118] ,
    \top_I.branch[11].l_um_iw[117] ,
    \top_I.branch[11].l_um_iw[116] ,
    \top_I.branch[11].l_um_iw[115] ,
    \top_I.branch[11].l_um_iw[114] ,
    \top_I.branch[11].l_um_iw[113] ,
    \top_I.branch[11].l_um_iw[112] ,
    \top_I.branch[11].l_um_iw[111] ,
    \top_I.branch[11].l_um_iw[110] ,
    \top_I.branch[11].l_um_iw[109] ,
    \top_I.branch[11].l_um_iw[108] ,
    \top_I.branch[11].l_um_iw[107] ,
    \top_I.branch[11].l_um_iw[106] ,
    \top_I.branch[11].l_um_iw[105] ,
    \top_I.branch[11].l_um_iw[104] ,
    \top_I.branch[11].l_um_iw[103] ,
    \top_I.branch[11].l_um_iw[102] ,
    \top_I.branch[11].l_um_iw[101] ,
    \top_I.branch[11].l_um_iw[100] ,
    \top_I.branch[11].l_um_iw[99] ,
    \top_I.branch[11].l_um_iw[98] ,
    \top_I.branch[11].l_um_iw[97] ,
    \top_I.branch[11].l_um_iw[96] ,
    \top_I.branch[11].l_um_iw[95] ,
    \top_I.branch[11].l_um_iw[94] ,
    \top_I.branch[11].l_um_iw[93] ,
    \top_I.branch[11].l_um_iw[92] ,
    \top_I.branch[11].l_um_iw[91] ,
    \top_I.branch[11].l_um_iw[90] ,
    \top_I.branch[11].l_um_iw[89] ,
    \top_I.branch[11].l_um_iw[88] ,
    \top_I.branch[11].l_um_iw[87] ,
    \top_I.branch[11].l_um_iw[86] ,
    \top_I.branch[11].l_um_iw[85] ,
    \top_I.branch[11].l_um_iw[84] ,
    \top_I.branch[11].l_um_iw[83] ,
    \top_I.branch[11].l_um_iw[82] ,
    \top_I.branch[11].l_um_iw[81] ,
    \top_I.branch[11].l_um_iw[80] ,
    \top_I.branch[11].l_um_iw[79] ,
    \top_I.branch[11].l_um_iw[78] ,
    \top_I.branch[11].l_um_iw[77] ,
    \top_I.branch[11].l_um_iw[76] ,
    \top_I.branch[11].l_um_iw[75] ,
    \top_I.branch[11].l_um_iw[74] ,
    \top_I.branch[11].l_um_iw[73] ,
    \top_I.branch[11].l_um_iw[72] ,
    \top_I.branch[11].l_um_iw[71] ,
    \top_I.branch[11].l_um_iw[70] ,
    \top_I.branch[11].l_um_iw[69] ,
    \top_I.branch[11].l_um_iw[68] ,
    \top_I.branch[11].l_um_iw[67] ,
    \top_I.branch[11].l_um_iw[66] ,
    \top_I.branch[11].l_um_iw[65] ,
    \top_I.branch[11].l_um_iw[64] ,
    \top_I.branch[11].l_um_iw[63] ,
    \top_I.branch[11].l_um_iw[62] ,
    \top_I.branch[11].l_um_iw[61] ,
    \top_I.branch[11].l_um_iw[60] ,
    \top_I.branch[11].l_um_iw[59] ,
    \top_I.branch[11].l_um_iw[58] ,
    \top_I.branch[11].l_um_iw[57] ,
    \top_I.branch[11].l_um_iw[56] ,
    \top_I.branch[11].l_um_iw[55] ,
    \top_I.branch[11].l_um_iw[54] ,
    \top_I.branch[11].l_um_iw[53] ,
    \top_I.branch[11].l_um_iw[52] ,
    \top_I.branch[11].l_um_iw[51] ,
    \top_I.branch[11].l_um_iw[50] ,
    \top_I.branch[11].l_um_iw[49] ,
    \top_I.branch[11].l_um_iw[48] ,
    \top_I.branch[11].l_um_iw[47] ,
    \top_I.branch[11].l_um_iw[46] ,
    \top_I.branch[11].l_um_iw[45] ,
    \top_I.branch[11].l_um_iw[44] ,
    \top_I.branch[11].l_um_iw[43] ,
    \top_I.branch[11].l_um_iw[42] ,
    \top_I.branch[11].l_um_iw[41] ,
    \top_I.branch[11].l_um_iw[40] ,
    \top_I.branch[11].l_um_iw[39] ,
    \top_I.branch[11].l_um_iw[38] ,
    \top_I.branch[11].l_um_iw[37] ,
    \top_I.branch[11].l_um_iw[36] ,
    \top_I.branch[11].l_um_iw[35] ,
    \top_I.branch[11].l_um_iw[34] ,
    \top_I.branch[11].l_um_iw[33] ,
    \top_I.branch[11].l_um_iw[32] ,
    \top_I.branch[11].l_um_iw[31] ,
    \top_I.branch[11].l_um_iw[30] ,
    \top_I.branch[11].l_um_iw[29] ,
    \top_I.branch[11].l_um_iw[28] ,
    \top_I.branch[11].l_um_iw[27] ,
    \top_I.branch[11].l_um_iw[26] ,
    \top_I.branch[11].l_um_iw[25] ,
    \top_I.branch[11].l_um_iw[24] ,
    \top_I.branch[11].l_um_iw[23] ,
    \top_I.branch[11].l_um_iw[22] ,
    \top_I.branch[11].l_um_iw[21] ,
    \top_I.branch[11].l_um_iw[20] ,
    \top_I.branch[11].l_um_iw[19] ,
    \top_I.branch[11].l_um_iw[18] ,
    \top_I.branch[11].l_um_iw[17] ,
    \top_I.branch[11].l_um_iw[16] ,
    \top_I.branch[11].l_um_iw[15] ,
    \top_I.branch[11].l_um_iw[14] ,
    \top_I.branch[11].l_um_iw[13] ,
    \top_I.branch[11].l_um_iw[12] ,
    \top_I.branch[11].l_um_iw[11] ,
    \top_I.branch[11].l_um_iw[10] ,
    \top_I.branch[11].l_um_iw[9] ,
    \top_I.branch[11].l_um_iw[8] ,
    \top_I.branch[11].l_um_iw[7] ,
    \top_I.branch[11].l_um_iw[6] ,
    \top_I.branch[11].l_um_iw[5] ,
    \top_I.branch[11].l_um_iw[4] ,
    \top_I.branch[11].l_um_iw[3] ,
    \top_I.branch[11].l_um_iw[2] ,
    \top_I.branch[11].l_um_iw[1] ,
    \top_I.branch[11].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[1] ,
    \top_I.branch[11].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[15] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[14] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[13] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[12] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[11] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[10] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[9] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[8] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[7] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[6] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[5] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[4] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[3] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].l_um_k_zero[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[11].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] ,
    \top_I.branch[11].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[12].col_um[0].um_bot_I.block_12_0.tt_um_I  (.clk(\top_I.branch[12].l_um_iw[0] ),
    .ena(\top_I.branch[12].l_um_ena[0] ),
    .rst_n(\top_I.branch[12].l_um_iw[1] ),
    .ui_in({\top_I.branch[12].l_um_iw[9] ,
    \top_I.branch[12].l_um_iw[8] ,
    \top_I.branch[12].l_um_iw[7] ,
    \top_I.branch[12].l_um_iw[6] ,
    \top_I.branch[12].l_um_iw[5] ,
    \top_I.branch[12].l_um_iw[4] ,
    \top_I.branch[12].l_um_iw[3] ,
    \top_I.branch[12].l_um_iw[2] }),
    .uio_in({\top_I.branch[12].l_um_iw[17] ,
    \top_I.branch[12].l_um_iw[16] ,
    \top_I.branch[12].l_um_iw[15] ,
    \top_I.branch[12].l_um_iw[14] ,
    \top_I.branch[12].l_um_iw[13] ,
    \top_I.branch[12].l_um_iw[12] ,
    \top_I.branch[12].l_um_iw[11] ,
    \top_I.branch[12].l_um_iw[10] }),
    .uio_oe({\top_I.branch[12].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[12].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[12].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[12].mux_I  (.k_one(\top_I.branch[12].l_k_one ),
    .k_zero(\top_I.branch[12].l_k_zero ),
    .addr({\top_I.branch[12].l_k_zero ,
    \top_I.branch[12].l_k_one ,
    \top_I.branch[12].l_k_one ,
    \top_I.branch[12].l_k_zero ,
    \top_I.branch[12].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[12].l_um_ena[15] ,
    \top_I.branch[12].l_um_ena[14] ,
    \top_I.branch[12].l_um_ena[13] ,
    \top_I.branch[12].l_um_ena[12] ,
    \top_I.branch[12].l_um_ena[11] ,
    \top_I.branch[12].l_um_ena[10] ,
    \top_I.branch[12].l_um_ena[9] ,
    \top_I.branch[12].l_um_ena[8] ,
    \top_I.branch[12].l_um_ena[7] ,
    \top_I.branch[12].l_um_ena[6] ,
    \top_I.branch[12].l_um_ena[5] ,
    \top_I.branch[12].l_um_ena[4] ,
    \top_I.branch[12].l_um_ena[3] ,
    \top_I.branch[12].l_um_ena[2] ,
    \top_I.branch[12].l_um_ena[1] ,
    \top_I.branch[12].l_um_ena[0] }),
    .um_iw({\top_I.branch[12].l_um_iw[287] ,
    \top_I.branch[12].l_um_iw[286] ,
    \top_I.branch[12].l_um_iw[285] ,
    \top_I.branch[12].l_um_iw[284] ,
    \top_I.branch[12].l_um_iw[283] ,
    \top_I.branch[12].l_um_iw[282] ,
    \top_I.branch[12].l_um_iw[281] ,
    \top_I.branch[12].l_um_iw[280] ,
    \top_I.branch[12].l_um_iw[279] ,
    \top_I.branch[12].l_um_iw[278] ,
    \top_I.branch[12].l_um_iw[277] ,
    \top_I.branch[12].l_um_iw[276] ,
    \top_I.branch[12].l_um_iw[275] ,
    \top_I.branch[12].l_um_iw[274] ,
    \top_I.branch[12].l_um_iw[273] ,
    \top_I.branch[12].l_um_iw[272] ,
    \top_I.branch[12].l_um_iw[271] ,
    \top_I.branch[12].l_um_iw[270] ,
    \top_I.branch[12].l_um_iw[269] ,
    \top_I.branch[12].l_um_iw[268] ,
    \top_I.branch[12].l_um_iw[267] ,
    \top_I.branch[12].l_um_iw[266] ,
    \top_I.branch[12].l_um_iw[265] ,
    \top_I.branch[12].l_um_iw[264] ,
    \top_I.branch[12].l_um_iw[263] ,
    \top_I.branch[12].l_um_iw[262] ,
    \top_I.branch[12].l_um_iw[261] ,
    \top_I.branch[12].l_um_iw[260] ,
    \top_I.branch[12].l_um_iw[259] ,
    \top_I.branch[12].l_um_iw[258] ,
    \top_I.branch[12].l_um_iw[257] ,
    \top_I.branch[12].l_um_iw[256] ,
    \top_I.branch[12].l_um_iw[255] ,
    \top_I.branch[12].l_um_iw[254] ,
    \top_I.branch[12].l_um_iw[253] ,
    \top_I.branch[12].l_um_iw[252] ,
    \top_I.branch[12].l_um_iw[251] ,
    \top_I.branch[12].l_um_iw[250] ,
    \top_I.branch[12].l_um_iw[249] ,
    \top_I.branch[12].l_um_iw[248] ,
    \top_I.branch[12].l_um_iw[247] ,
    \top_I.branch[12].l_um_iw[246] ,
    \top_I.branch[12].l_um_iw[245] ,
    \top_I.branch[12].l_um_iw[244] ,
    \top_I.branch[12].l_um_iw[243] ,
    \top_I.branch[12].l_um_iw[242] ,
    \top_I.branch[12].l_um_iw[241] ,
    \top_I.branch[12].l_um_iw[240] ,
    \top_I.branch[12].l_um_iw[239] ,
    \top_I.branch[12].l_um_iw[238] ,
    \top_I.branch[12].l_um_iw[237] ,
    \top_I.branch[12].l_um_iw[236] ,
    \top_I.branch[12].l_um_iw[235] ,
    \top_I.branch[12].l_um_iw[234] ,
    \top_I.branch[12].l_um_iw[233] ,
    \top_I.branch[12].l_um_iw[232] ,
    \top_I.branch[12].l_um_iw[231] ,
    \top_I.branch[12].l_um_iw[230] ,
    \top_I.branch[12].l_um_iw[229] ,
    \top_I.branch[12].l_um_iw[228] ,
    \top_I.branch[12].l_um_iw[227] ,
    \top_I.branch[12].l_um_iw[226] ,
    \top_I.branch[12].l_um_iw[225] ,
    \top_I.branch[12].l_um_iw[224] ,
    \top_I.branch[12].l_um_iw[223] ,
    \top_I.branch[12].l_um_iw[222] ,
    \top_I.branch[12].l_um_iw[221] ,
    \top_I.branch[12].l_um_iw[220] ,
    \top_I.branch[12].l_um_iw[219] ,
    \top_I.branch[12].l_um_iw[218] ,
    \top_I.branch[12].l_um_iw[217] ,
    \top_I.branch[12].l_um_iw[216] ,
    \top_I.branch[12].l_um_iw[215] ,
    \top_I.branch[12].l_um_iw[214] ,
    \top_I.branch[12].l_um_iw[213] ,
    \top_I.branch[12].l_um_iw[212] ,
    \top_I.branch[12].l_um_iw[211] ,
    \top_I.branch[12].l_um_iw[210] ,
    \top_I.branch[12].l_um_iw[209] ,
    \top_I.branch[12].l_um_iw[208] ,
    \top_I.branch[12].l_um_iw[207] ,
    \top_I.branch[12].l_um_iw[206] ,
    \top_I.branch[12].l_um_iw[205] ,
    \top_I.branch[12].l_um_iw[204] ,
    \top_I.branch[12].l_um_iw[203] ,
    \top_I.branch[12].l_um_iw[202] ,
    \top_I.branch[12].l_um_iw[201] ,
    \top_I.branch[12].l_um_iw[200] ,
    \top_I.branch[12].l_um_iw[199] ,
    \top_I.branch[12].l_um_iw[198] ,
    \top_I.branch[12].l_um_iw[197] ,
    \top_I.branch[12].l_um_iw[196] ,
    \top_I.branch[12].l_um_iw[195] ,
    \top_I.branch[12].l_um_iw[194] ,
    \top_I.branch[12].l_um_iw[193] ,
    \top_I.branch[12].l_um_iw[192] ,
    \top_I.branch[12].l_um_iw[191] ,
    \top_I.branch[12].l_um_iw[190] ,
    \top_I.branch[12].l_um_iw[189] ,
    \top_I.branch[12].l_um_iw[188] ,
    \top_I.branch[12].l_um_iw[187] ,
    \top_I.branch[12].l_um_iw[186] ,
    \top_I.branch[12].l_um_iw[185] ,
    \top_I.branch[12].l_um_iw[184] ,
    \top_I.branch[12].l_um_iw[183] ,
    \top_I.branch[12].l_um_iw[182] ,
    \top_I.branch[12].l_um_iw[181] ,
    \top_I.branch[12].l_um_iw[180] ,
    \top_I.branch[12].l_um_iw[179] ,
    \top_I.branch[12].l_um_iw[178] ,
    \top_I.branch[12].l_um_iw[177] ,
    \top_I.branch[12].l_um_iw[176] ,
    \top_I.branch[12].l_um_iw[175] ,
    \top_I.branch[12].l_um_iw[174] ,
    \top_I.branch[12].l_um_iw[173] ,
    \top_I.branch[12].l_um_iw[172] ,
    \top_I.branch[12].l_um_iw[171] ,
    \top_I.branch[12].l_um_iw[170] ,
    \top_I.branch[12].l_um_iw[169] ,
    \top_I.branch[12].l_um_iw[168] ,
    \top_I.branch[12].l_um_iw[167] ,
    \top_I.branch[12].l_um_iw[166] ,
    \top_I.branch[12].l_um_iw[165] ,
    \top_I.branch[12].l_um_iw[164] ,
    \top_I.branch[12].l_um_iw[163] ,
    \top_I.branch[12].l_um_iw[162] ,
    \top_I.branch[12].l_um_iw[161] ,
    \top_I.branch[12].l_um_iw[160] ,
    \top_I.branch[12].l_um_iw[159] ,
    \top_I.branch[12].l_um_iw[158] ,
    \top_I.branch[12].l_um_iw[157] ,
    \top_I.branch[12].l_um_iw[156] ,
    \top_I.branch[12].l_um_iw[155] ,
    \top_I.branch[12].l_um_iw[154] ,
    \top_I.branch[12].l_um_iw[153] ,
    \top_I.branch[12].l_um_iw[152] ,
    \top_I.branch[12].l_um_iw[151] ,
    \top_I.branch[12].l_um_iw[150] ,
    \top_I.branch[12].l_um_iw[149] ,
    \top_I.branch[12].l_um_iw[148] ,
    \top_I.branch[12].l_um_iw[147] ,
    \top_I.branch[12].l_um_iw[146] ,
    \top_I.branch[12].l_um_iw[145] ,
    \top_I.branch[12].l_um_iw[144] ,
    \top_I.branch[12].l_um_iw[143] ,
    \top_I.branch[12].l_um_iw[142] ,
    \top_I.branch[12].l_um_iw[141] ,
    \top_I.branch[12].l_um_iw[140] ,
    \top_I.branch[12].l_um_iw[139] ,
    \top_I.branch[12].l_um_iw[138] ,
    \top_I.branch[12].l_um_iw[137] ,
    \top_I.branch[12].l_um_iw[136] ,
    \top_I.branch[12].l_um_iw[135] ,
    \top_I.branch[12].l_um_iw[134] ,
    \top_I.branch[12].l_um_iw[133] ,
    \top_I.branch[12].l_um_iw[132] ,
    \top_I.branch[12].l_um_iw[131] ,
    \top_I.branch[12].l_um_iw[130] ,
    \top_I.branch[12].l_um_iw[129] ,
    \top_I.branch[12].l_um_iw[128] ,
    \top_I.branch[12].l_um_iw[127] ,
    \top_I.branch[12].l_um_iw[126] ,
    \top_I.branch[12].l_um_iw[125] ,
    \top_I.branch[12].l_um_iw[124] ,
    \top_I.branch[12].l_um_iw[123] ,
    \top_I.branch[12].l_um_iw[122] ,
    \top_I.branch[12].l_um_iw[121] ,
    \top_I.branch[12].l_um_iw[120] ,
    \top_I.branch[12].l_um_iw[119] ,
    \top_I.branch[12].l_um_iw[118] ,
    \top_I.branch[12].l_um_iw[117] ,
    \top_I.branch[12].l_um_iw[116] ,
    \top_I.branch[12].l_um_iw[115] ,
    \top_I.branch[12].l_um_iw[114] ,
    \top_I.branch[12].l_um_iw[113] ,
    \top_I.branch[12].l_um_iw[112] ,
    \top_I.branch[12].l_um_iw[111] ,
    \top_I.branch[12].l_um_iw[110] ,
    \top_I.branch[12].l_um_iw[109] ,
    \top_I.branch[12].l_um_iw[108] ,
    \top_I.branch[12].l_um_iw[107] ,
    \top_I.branch[12].l_um_iw[106] ,
    \top_I.branch[12].l_um_iw[105] ,
    \top_I.branch[12].l_um_iw[104] ,
    \top_I.branch[12].l_um_iw[103] ,
    \top_I.branch[12].l_um_iw[102] ,
    \top_I.branch[12].l_um_iw[101] ,
    \top_I.branch[12].l_um_iw[100] ,
    \top_I.branch[12].l_um_iw[99] ,
    \top_I.branch[12].l_um_iw[98] ,
    \top_I.branch[12].l_um_iw[97] ,
    \top_I.branch[12].l_um_iw[96] ,
    \top_I.branch[12].l_um_iw[95] ,
    \top_I.branch[12].l_um_iw[94] ,
    \top_I.branch[12].l_um_iw[93] ,
    \top_I.branch[12].l_um_iw[92] ,
    \top_I.branch[12].l_um_iw[91] ,
    \top_I.branch[12].l_um_iw[90] ,
    \top_I.branch[12].l_um_iw[89] ,
    \top_I.branch[12].l_um_iw[88] ,
    \top_I.branch[12].l_um_iw[87] ,
    \top_I.branch[12].l_um_iw[86] ,
    \top_I.branch[12].l_um_iw[85] ,
    \top_I.branch[12].l_um_iw[84] ,
    \top_I.branch[12].l_um_iw[83] ,
    \top_I.branch[12].l_um_iw[82] ,
    \top_I.branch[12].l_um_iw[81] ,
    \top_I.branch[12].l_um_iw[80] ,
    \top_I.branch[12].l_um_iw[79] ,
    \top_I.branch[12].l_um_iw[78] ,
    \top_I.branch[12].l_um_iw[77] ,
    \top_I.branch[12].l_um_iw[76] ,
    \top_I.branch[12].l_um_iw[75] ,
    \top_I.branch[12].l_um_iw[74] ,
    \top_I.branch[12].l_um_iw[73] ,
    \top_I.branch[12].l_um_iw[72] ,
    \top_I.branch[12].l_um_iw[71] ,
    \top_I.branch[12].l_um_iw[70] ,
    \top_I.branch[12].l_um_iw[69] ,
    \top_I.branch[12].l_um_iw[68] ,
    \top_I.branch[12].l_um_iw[67] ,
    \top_I.branch[12].l_um_iw[66] ,
    \top_I.branch[12].l_um_iw[65] ,
    \top_I.branch[12].l_um_iw[64] ,
    \top_I.branch[12].l_um_iw[63] ,
    \top_I.branch[12].l_um_iw[62] ,
    \top_I.branch[12].l_um_iw[61] ,
    \top_I.branch[12].l_um_iw[60] ,
    \top_I.branch[12].l_um_iw[59] ,
    \top_I.branch[12].l_um_iw[58] ,
    \top_I.branch[12].l_um_iw[57] ,
    \top_I.branch[12].l_um_iw[56] ,
    \top_I.branch[12].l_um_iw[55] ,
    \top_I.branch[12].l_um_iw[54] ,
    \top_I.branch[12].l_um_iw[53] ,
    \top_I.branch[12].l_um_iw[52] ,
    \top_I.branch[12].l_um_iw[51] ,
    \top_I.branch[12].l_um_iw[50] ,
    \top_I.branch[12].l_um_iw[49] ,
    \top_I.branch[12].l_um_iw[48] ,
    \top_I.branch[12].l_um_iw[47] ,
    \top_I.branch[12].l_um_iw[46] ,
    \top_I.branch[12].l_um_iw[45] ,
    \top_I.branch[12].l_um_iw[44] ,
    \top_I.branch[12].l_um_iw[43] ,
    \top_I.branch[12].l_um_iw[42] ,
    \top_I.branch[12].l_um_iw[41] ,
    \top_I.branch[12].l_um_iw[40] ,
    \top_I.branch[12].l_um_iw[39] ,
    \top_I.branch[12].l_um_iw[38] ,
    \top_I.branch[12].l_um_iw[37] ,
    \top_I.branch[12].l_um_iw[36] ,
    \top_I.branch[12].l_um_iw[35] ,
    \top_I.branch[12].l_um_iw[34] ,
    \top_I.branch[12].l_um_iw[33] ,
    \top_I.branch[12].l_um_iw[32] ,
    \top_I.branch[12].l_um_iw[31] ,
    \top_I.branch[12].l_um_iw[30] ,
    \top_I.branch[12].l_um_iw[29] ,
    \top_I.branch[12].l_um_iw[28] ,
    \top_I.branch[12].l_um_iw[27] ,
    \top_I.branch[12].l_um_iw[26] ,
    \top_I.branch[12].l_um_iw[25] ,
    \top_I.branch[12].l_um_iw[24] ,
    \top_I.branch[12].l_um_iw[23] ,
    \top_I.branch[12].l_um_iw[22] ,
    \top_I.branch[12].l_um_iw[21] ,
    \top_I.branch[12].l_um_iw[20] ,
    \top_I.branch[12].l_um_iw[19] ,
    \top_I.branch[12].l_um_iw[18] ,
    \top_I.branch[12].l_um_iw[17] ,
    \top_I.branch[12].l_um_iw[16] ,
    \top_I.branch[12].l_um_iw[15] ,
    \top_I.branch[12].l_um_iw[14] ,
    \top_I.branch[12].l_um_iw[13] ,
    \top_I.branch[12].l_um_iw[12] ,
    \top_I.branch[12].l_um_iw[11] ,
    \top_I.branch[12].l_um_iw[10] ,
    \top_I.branch[12].l_um_iw[9] ,
    \top_I.branch[12].l_um_iw[8] ,
    \top_I.branch[12].l_um_iw[7] ,
    \top_I.branch[12].l_um_iw[6] ,
    \top_I.branch[12].l_um_iw[5] ,
    \top_I.branch[12].l_um_iw[4] ,
    \top_I.branch[12].l_um_iw[3] ,
    \top_I.branch[12].l_um_iw[2] ,
    \top_I.branch[12].l_um_iw[1] ,
    \top_I.branch[12].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[15] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[14] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[13] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[12] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[11] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[10] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[9] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[8] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[7] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[6] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[5] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[4] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[3] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[2] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].l_um_k_zero[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[12].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[13].col_um[0].um_bot_I.block_12_16.tt_um_I  (.clk(\top_I.branch[13].l_um_iw[0] ),
    .ena(\top_I.branch[13].l_um_ena[0] ),
    .rst_n(\top_I.branch[13].l_um_iw[1] ),
    .ui_in({\top_I.branch[13].l_um_iw[9] ,
    \top_I.branch[13].l_um_iw[8] ,
    \top_I.branch[13].l_um_iw[7] ,
    \top_I.branch[13].l_um_iw[6] ,
    \top_I.branch[13].l_um_iw[5] ,
    \top_I.branch[13].l_um_iw[4] ,
    \top_I.branch[13].l_um_iw[3] ,
    \top_I.branch[13].l_um_iw[2] }),
    .uio_in({\top_I.branch[13].l_um_iw[17] ,
    \top_I.branch[13].l_um_iw[16] ,
    \top_I.branch[13].l_um_iw[15] ,
    \top_I.branch[13].l_um_iw[14] ,
    \top_I.branch[13].l_um_iw[13] ,
    \top_I.branch[13].l_um_iw[12] ,
    \top_I.branch[13].l_um_iw[11] ,
    \top_I.branch[13].l_um_iw[10] }),
    .uio_oe({\top_I.branch[13].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[13].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[13].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[13].mux_I  (.k_one(\top_I.branch[13].l_k_one ),
    .k_zero(\top_I.branch[13].l_k_zero ),
    .addr({\top_I.branch[13].l_k_zero ,
    \top_I.branch[13].l_k_one ,
    \top_I.branch[13].l_k_one ,
    \top_I.branch[13].l_k_zero ,
    \top_I.branch[13].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[13].l_um_ena[15] ,
    \top_I.branch[13].l_um_ena[14] ,
    \top_I.branch[13].l_um_ena[13] ,
    \top_I.branch[13].l_um_ena[12] ,
    \top_I.branch[13].l_um_ena[11] ,
    \top_I.branch[13].l_um_ena[10] ,
    \top_I.branch[13].l_um_ena[9] ,
    \top_I.branch[13].l_um_ena[8] ,
    \top_I.branch[13].l_um_ena[7] ,
    \top_I.branch[13].l_um_ena[6] ,
    \top_I.branch[13].l_um_ena[5] ,
    \top_I.branch[13].l_um_ena[4] ,
    \top_I.branch[13].l_um_ena[3] ,
    \top_I.branch[13].l_um_ena[2] ,
    \top_I.branch[13].l_um_ena[1] ,
    \top_I.branch[13].l_um_ena[0] }),
    .um_iw({\top_I.branch[13].l_um_iw[287] ,
    \top_I.branch[13].l_um_iw[286] ,
    \top_I.branch[13].l_um_iw[285] ,
    \top_I.branch[13].l_um_iw[284] ,
    \top_I.branch[13].l_um_iw[283] ,
    \top_I.branch[13].l_um_iw[282] ,
    \top_I.branch[13].l_um_iw[281] ,
    \top_I.branch[13].l_um_iw[280] ,
    \top_I.branch[13].l_um_iw[279] ,
    \top_I.branch[13].l_um_iw[278] ,
    \top_I.branch[13].l_um_iw[277] ,
    \top_I.branch[13].l_um_iw[276] ,
    \top_I.branch[13].l_um_iw[275] ,
    \top_I.branch[13].l_um_iw[274] ,
    \top_I.branch[13].l_um_iw[273] ,
    \top_I.branch[13].l_um_iw[272] ,
    \top_I.branch[13].l_um_iw[271] ,
    \top_I.branch[13].l_um_iw[270] ,
    \top_I.branch[13].l_um_iw[269] ,
    \top_I.branch[13].l_um_iw[268] ,
    \top_I.branch[13].l_um_iw[267] ,
    \top_I.branch[13].l_um_iw[266] ,
    \top_I.branch[13].l_um_iw[265] ,
    \top_I.branch[13].l_um_iw[264] ,
    \top_I.branch[13].l_um_iw[263] ,
    \top_I.branch[13].l_um_iw[262] ,
    \top_I.branch[13].l_um_iw[261] ,
    \top_I.branch[13].l_um_iw[260] ,
    \top_I.branch[13].l_um_iw[259] ,
    \top_I.branch[13].l_um_iw[258] ,
    \top_I.branch[13].l_um_iw[257] ,
    \top_I.branch[13].l_um_iw[256] ,
    \top_I.branch[13].l_um_iw[255] ,
    \top_I.branch[13].l_um_iw[254] ,
    \top_I.branch[13].l_um_iw[253] ,
    \top_I.branch[13].l_um_iw[252] ,
    \top_I.branch[13].l_um_iw[251] ,
    \top_I.branch[13].l_um_iw[250] ,
    \top_I.branch[13].l_um_iw[249] ,
    \top_I.branch[13].l_um_iw[248] ,
    \top_I.branch[13].l_um_iw[247] ,
    \top_I.branch[13].l_um_iw[246] ,
    \top_I.branch[13].l_um_iw[245] ,
    \top_I.branch[13].l_um_iw[244] ,
    \top_I.branch[13].l_um_iw[243] ,
    \top_I.branch[13].l_um_iw[242] ,
    \top_I.branch[13].l_um_iw[241] ,
    \top_I.branch[13].l_um_iw[240] ,
    \top_I.branch[13].l_um_iw[239] ,
    \top_I.branch[13].l_um_iw[238] ,
    \top_I.branch[13].l_um_iw[237] ,
    \top_I.branch[13].l_um_iw[236] ,
    \top_I.branch[13].l_um_iw[235] ,
    \top_I.branch[13].l_um_iw[234] ,
    \top_I.branch[13].l_um_iw[233] ,
    \top_I.branch[13].l_um_iw[232] ,
    \top_I.branch[13].l_um_iw[231] ,
    \top_I.branch[13].l_um_iw[230] ,
    \top_I.branch[13].l_um_iw[229] ,
    \top_I.branch[13].l_um_iw[228] ,
    \top_I.branch[13].l_um_iw[227] ,
    \top_I.branch[13].l_um_iw[226] ,
    \top_I.branch[13].l_um_iw[225] ,
    \top_I.branch[13].l_um_iw[224] ,
    \top_I.branch[13].l_um_iw[223] ,
    \top_I.branch[13].l_um_iw[222] ,
    \top_I.branch[13].l_um_iw[221] ,
    \top_I.branch[13].l_um_iw[220] ,
    \top_I.branch[13].l_um_iw[219] ,
    \top_I.branch[13].l_um_iw[218] ,
    \top_I.branch[13].l_um_iw[217] ,
    \top_I.branch[13].l_um_iw[216] ,
    \top_I.branch[13].l_um_iw[215] ,
    \top_I.branch[13].l_um_iw[214] ,
    \top_I.branch[13].l_um_iw[213] ,
    \top_I.branch[13].l_um_iw[212] ,
    \top_I.branch[13].l_um_iw[211] ,
    \top_I.branch[13].l_um_iw[210] ,
    \top_I.branch[13].l_um_iw[209] ,
    \top_I.branch[13].l_um_iw[208] ,
    \top_I.branch[13].l_um_iw[207] ,
    \top_I.branch[13].l_um_iw[206] ,
    \top_I.branch[13].l_um_iw[205] ,
    \top_I.branch[13].l_um_iw[204] ,
    \top_I.branch[13].l_um_iw[203] ,
    \top_I.branch[13].l_um_iw[202] ,
    \top_I.branch[13].l_um_iw[201] ,
    \top_I.branch[13].l_um_iw[200] ,
    \top_I.branch[13].l_um_iw[199] ,
    \top_I.branch[13].l_um_iw[198] ,
    \top_I.branch[13].l_um_iw[197] ,
    \top_I.branch[13].l_um_iw[196] ,
    \top_I.branch[13].l_um_iw[195] ,
    \top_I.branch[13].l_um_iw[194] ,
    \top_I.branch[13].l_um_iw[193] ,
    \top_I.branch[13].l_um_iw[192] ,
    \top_I.branch[13].l_um_iw[191] ,
    \top_I.branch[13].l_um_iw[190] ,
    \top_I.branch[13].l_um_iw[189] ,
    \top_I.branch[13].l_um_iw[188] ,
    \top_I.branch[13].l_um_iw[187] ,
    \top_I.branch[13].l_um_iw[186] ,
    \top_I.branch[13].l_um_iw[185] ,
    \top_I.branch[13].l_um_iw[184] ,
    \top_I.branch[13].l_um_iw[183] ,
    \top_I.branch[13].l_um_iw[182] ,
    \top_I.branch[13].l_um_iw[181] ,
    \top_I.branch[13].l_um_iw[180] ,
    \top_I.branch[13].l_um_iw[179] ,
    \top_I.branch[13].l_um_iw[178] ,
    \top_I.branch[13].l_um_iw[177] ,
    \top_I.branch[13].l_um_iw[176] ,
    \top_I.branch[13].l_um_iw[175] ,
    \top_I.branch[13].l_um_iw[174] ,
    \top_I.branch[13].l_um_iw[173] ,
    \top_I.branch[13].l_um_iw[172] ,
    \top_I.branch[13].l_um_iw[171] ,
    \top_I.branch[13].l_um_iw[170] ,
    \top_I.branch[13].l_um_iw[169] ,
    \top_I.branch[13].l_um_iw[168] ,
    \top_I.branch[13].l_um_iw[167] ,
    \top_I.branch[13].l_um_iw[166] ,
    \top_I.branch[13].l_um_iw[165] ,
    \top_I.branch[13].l_um_iw[164] ,
    \top_I.branch[13].l_um_iw[163] ,
    \top_I.branch[13].l_um_iw[162] ,
    \top_I.branch[13].l_um_iw[161] ,
    \top_I.branch[13].l_um_iw[160] ,
    \top_I.branch[13].l_um_iw[159] ,
    \top_I.branch[13].l_um_iw[158] ,
    \top_I.branch[13].l_um_iw[157] ,
    \top_I.branch[13].l_um_iw[156] ,
    \top_I.branch[13].l_um_iw[155] ,
    \top_I.branch[13].l_um_iw[154] ,
    \top_I.branch[13].l_um_iw[153] ,
    \top_I.branch[13].l_um_iw[152] ,
    \top_I.branch[13].l_um_iw[151] ,
    \top_I.branch[13].l_um_iw[150] ,
    \top_I.branch[13].l_um_iw[149] ,
    \top_I.branch[13].l_um_iw[148] ,
    \top_I.branch[13].l_um_iw[147] ,
    \top_I.branch[13].l_um_iw[146] ,
    \top_I.branch[13].l_um_iw[145] ,
    \top_I.branch[13].l_um_iw[144] ,
    \top_I.branch[13].l_um_iw[143] ,
    \top_I.branch[13].l_um_iw[142] ,
    \top_I.branch[13].l_um_iw[141] ,
    \top_I.branch[13].l_um_iw[140] ,
    \top_I.branch[13].l_um_iw[139] ,
    \top_I.branch[13].l_um_iw[138] ,
    \top_I.branch[13].l_um_iw[137] ,
    \top_I.branch[13].l_um_iw[136] ,
    \top_I.branch[13].l_um_iw[135] ,
    \top_I.branch[13].l_um_iw[134] ,
    \top_I.branch[13].l_um_iw[133] ,
    \top_I.branch[13].l_um_iw[132] ,
    \top_I.branch[13].l_um_iw[131] ,
    \top_I.branch[13].l_um_iw[130] ,
    \top_I.branch[13].l_um_iw[129] ,
    \top_I.branch[13].l_um_iw[128] ,
    \top_I.branch[13].l_um_iw[127] ,
    \top_I.branch[13].l_um_iw[126] ,
    \top_I.branch[13].l_um_iw[125] ,
    \top_I.branch[13].l_um_iw[124] ,
    \top_I.branch[13].l_um_iw[123] ,
    \top_I.branch[13].l_um_iw[122] ,
    \top_I.branch[13].l_um_iw[121] ,
    \top_I.branch[13].l_um_iw[120] ,
    \top_I.branch[13].l_um_iw[119] ,
    \top_I.branch[13].l_um_iw[118] ,
    \top_I.branch[13].l_um_iw[117] ,
    \top_I.branch[13].l_um_iw[116] ,
    \top_I.branch[13].l_um_iw[115] ,
    \top_I.branch[13].l_um_iw[114] ,
    \top_I.branch[13].l_um_iw[113] ,
    \top_I.branch[13].l_um_iw[112] ,
    \top_I.branch[13].l_um_iw[111] ,
    \top_I.branch[13].l_um_iw[110] ,
    \top_I.branch[13].l_um_iw[109] ,
    \top_I.branch[13].l_um_iw[108] ,
    \top_I.branch[13].l_um_iw[107] ,
    \top_I.branch[13].l_um_iw[106] ,
    \top_I.branch[13].l_um_iw[105] ,
    \top_I.branch[13].l_um_iw[104] ,
    \top_I.branch[13].l_um_iw[103] ,
    \top_I.branch[13].l_um_iw[102] ,
    \top_I.branch[13].l_um_iw[101] ,
    \top_I.branch[13].l_um_iw[100] ,
    \top_I.branch[13].l_um_iw[99] ,
    \top_I.branch[13].l_um_iw[98] ,
    \top_I.branch[13].l_um_iw[97] ,
    \top_I.branch[13].l_um_iw[96] ,
    \top_I.branch[13].l_um_iw[95] ,
    \top_I.branch[13].l_um_iw[94] ,
    \top_I.branch[13].l_um_iw[93] ,
    \top_I.branch[13].l_um_iw[92] ,
    \top_I.branch[13].l_um_iw[91] ,
    \top_I.branch[13].l_um_iw[90] ,
    \top_I.branch[13].l_um_iw[89] ,
    \top_I.branch[13].l_um_iw[88] ,
    \top_I.branch[13].l_um_iw[87] ,
    \top_I.branch[13].l_um_iw[86] ,
    \top_I.branch[13].l_um_iw[85] ,
    \top_I.branch[13].l_um_iw[84] ,
    \top_I.branch[13].l_um_iw[83] ,
    \top_I.branch[13].l_um_iw[82] ,
    \top_I.branch[13].l_um_iw[81] ,
    \top_I.branch[13].l_um_iw[80] ,
    \top_I.branch[13].l_um_iw[79] ,
    \top_I.branch[13].l_um_iw[78] ,
    \top_I.branch[13].l_um_iw[77] ,
    \top_I.branch[13].l_um_iw[76] ,
    \top_I.branch[13].l_um_iw[75] ,
    \top_I.branch[13].l_um_iw[74] ,
    \top_I.branch[13].l_um_iw[73] ,
    \top_I.branch[13].l_um_iw[72] ,
    \top_I.branch[13].l_um_iw[71] ,
    \top_I.branch[13].l_um_iw[70] ,
    \top_I.branch[13].l_um_iw[69] ,
    \top_I.branch[13].l_um_iw[68] ,
    \top_I.branch[13].l_um_iw[67] ,
    \top_I.branch[13].l_um_iw[66] ,
    \top_I.branch[13].l_um_iw[65] ,
    \top_I.branch[13].l_um_iw[64] ,
    \top_I.branch[13].l_um_iw[63] ,
    \top_I.branch[13].l_um_iw[62] ,
    \top_I.branch[13].l_um_iw[61] ,
    \top_I.branch[13].l_um_iw[60] ,
    \top_I.branch[13].l_um_iw[59] ,
    \top_I.branch[13].l_um_iw[58] ,
    \top_I.branch[13].l_um_iw[57] ,
    \top_I.branch[13].l_um_iw[56] ,
    \top_I.branch[13].l_um_iw[55] ,
    \top_I.branch[13].l_um_iw[54] ,
    \top_I.branch[13].l_um_iw[53] ,
    \top_I.branch[13].l_um_iw[52] ,
    \top_I.branch[13].l_um_iw[51] ,
    \top_I.branch[13].l_um_iw[50] ,
    \top_I.branch[13].l_um_iw[49] ,
    \top_I.branch[13].l_um_iw[48] ,
    \top_I.branch[13].l_um_iw[47] ,
    \top_I.branch[13].l_um_iw[46] ,
    \top_I.branch[13].l_um_iw[45] ,
    \top_I.branch[13].l_um_iw[44] ,
    \top_I.branch[13].l_um_iw[43] ,
    \top_I.branch[13].l_um_iw[42] ,
    \top_I.branch[13].l_um_iw[41] ,
    \top_I.branch[13].l_um_iw[40] ,
    \top_I.branch[13].l_um_iw[39] ,
    \top_I.branch[13].l_um_iw[38] ,
    \top_I.branch[13].l_um_iw[37] ,
    \top_I.branch[13].l_um_iw[36] ,
    \top_I.branch[13].l_um_iw[35] ,
    \top_I.branch[13].l_um_iw[34] ,
    \top_I.branch[13].l_um_iw[33] ,
    \top_I.branch[13].l_um_iw[32] ,
    \top_I.branch[13].l_um_iw[31] ,
    \top_I.branch[13].l_um_iw[30] ,
    \top_I.branch[13].l_um_iw[29] ,
    \top_I.branch[13].l_um_iw[28] ,
    \top_I.branch[13].l_um_iw[27] ,
    \top_I.branch[13].l_um_iw[26] ,
    \top_I.branch[13].l_um_iw[25] ,
    \top_I.branch[13].l_um_iw[24] ,
    \top_I.branch[13].l_um_iw[23] ,
    \top_I.branch[13].l_um_iw[22] ,
    \top_I.branch[13].l_um_iw[21] ,
    \top_I.branch[13].l_um_iw[20] ,
    \top_I.branch[13].l_um_iw[19] ,
    \top_I.branch[13].l_um_iw[18] ,
    \top_I.branch[13].l_um_iw[17] ,
    \top_I.branch[13].l_um_iw[16] ,
    \top_I.branch[13].l_um_iw[15] ,
    \top_I.branch[13].l_um_iw[14] ,
    \top_I.branch[13].l_um_iw[13] ,
    \top_I.branch[13].l_um_iw[12] ,
    \top_I.branch[13].l_um_iw[11] ,
    \top_I.branch[13].l_um_iw[10] ,
    \top_I.branch[13].l_um_iw[9] ,
    \top_I.branch[13].l_um_iw[8] ,
    \top_I.branch[13].l_um_iw[7] ,
    \top_I.branch[13].l_um_iw[6] ,
    \top_I.branch[13].l_um_iw[5] ,
    \top_I.branch[13].l_um_iw[4] ,
    \top_I.branch[13].l_um_iw[3] ,
    \top_I.branch[13].l_um_iw[2] ,
    \top_I.branch[13].l_um_iw[1] ,
    \top_I.branch[13].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[15] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[14] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[13] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[12] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[11] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[10] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[9] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[8] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[7] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[6] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[5] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[4] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[3] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[2] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].l_um_k_zero[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[13].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[14].col_um[0].um_top_I.block_15_0.tt_um_I  (.clk(\top_I.branch[14].l_um_iw[18] ),
    .ena(\top_I.branch[14].l_um_ena[1] ),
    .rst_n(\top_I.branch[14].l_um_iw[19] ),
    .ui_in({\top_I.branch[14].l_um_iw[27] ,
    \top_I.branch[14].l_um_iw[26] ,
    \top_I.branch[14].l_um_iw[25] ,
    \top_I.branch[14].l_um_iw[24] ,
    \top_I.branch[14].l_um_iw[23] ,
    \top_I.branch[14].l_um_iw[22] ,
    \top_I.branch[14].l_um_iw[21] ,
    \top_I.branch[14].l_um_iw[20] }),
    .uio_in({\top_I.branch[14].l_um_iw[35] ,
    \top_I.branch[14].l_um_iw[34] ,
    \top_I.branch[14].l_um_iw[33] ,
    \top_I.branch[14].l_um_iw[32] ,
    \top_I.branch[14].l_um_iw[31] ,
    \top_I.branch[14].l_um_iw[30] ,
    \top_I.branch[14].l_um_iw[29] ,
    \top_I.branch[14].l_um_iw[28] }),
    .uio_oe({\top_I.branch[14].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[14].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[14].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[14].mux_I  (.k_one(\top_I.branch[14].l_k_one ),
    .k_zero(\top_I.branch[14].l_k_zero ),
    .addr({\top_I.branch[14].l_k_zero ,
    \top_I.branch[14].l_k_one ,
    \top_I.branch[14].l_k_one ,
    \top_I.branch[14].l_k_one ,
    \top_I.branch[14].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[14].l_um_ena[15] ,
    \top_I.branch[14].l_um_ena[14] ,
    \top_I.branch[14].l_um_ena[13] ,
    \top_I.branch[14].l_um_ena[12] ,
    \top_I.branch[14].l_um_ena[11] ,
    \top_I.branch[14].l_um_ena[10] ,
    \top_I.branch[14].l_um_ena[9] ,
    \top_I.branch[14].l_um_ena[8] ,
    \top_I.branch[14].l_um_ena[7] ,
    \top_I.branch[14].l_um_ena[6] ,
    \top_I.branch[14].l_um_ena[5] ,
    \top_I.branch[14].l_um_ena[4] ,
    \top_I.branch[14].l_um_ena[3] ,
    \top_I.branch[14].l_um_ena[2] ,
    \top_I.branch[14].l_um_ena[1] ,
    \top_I.branch[14].l_um_ena[0] }),
    .um_iw({\top_I.branch[14].l_um_iw[287] ,
    \top_I.branch[14].l_um_iw[286] ,
    \top_I.branch[14].l_um_iw[285] ,
    \top_I.branch[14].l_um_iw[284] ,
    \top_I.branch[14].l_um_iw[283] ,
    \top_I.branch[14].l_um_iw[282] ,
    \top_I.branch[14].l_um_iw[281] ,
    \top_I.branch[14].l_um_iw[280] ,
    \top_I.branch[14].l_um_iw[279] ,
    \top_I.branch[14].l_um_iw[278] ,
    \top_I.branch[14].l_um_iw[277] ,
    \top_I.branch[14].l_um_iw[276] ,
    \top_I.branch[14].l_um_iw[275] ,
    \top_I.branch[14].l_um_iw[274] ,
    \top_I.branch[14].l_um_iw[273] ,
    \top_I.branch[14].l_um_iw[272] ,
    \top_I.branch[14].l_um_iw[271] ,
    \top_I.branch[14].l_um_iw[270] ,
    \top_I.branch[14].l_um_iw[269] ,
    \top_I.branch[14].l_um_iw[268] ,
    \top_I.branch[14].l_um_iw[267] ,
    \top_I.branch[14].l_um_iw[266] ,
    \top_I.branch[14].l_um_iw[265] ,
    \top_I.branch[14].l_um_iw[264] ,
    \top_I.branch[14].l_um_iw[263] ,
    \top_I.branch[14].l_um_iw[262] ,
    \top_I.branch[14].l_um_iw[261] ,
    \top_I.branch[14].l_um_iw[260] ,
    \top_I.branch[14].l_um_iw[259] ,
    \top_I.branch[14].l_um_iw[258] ,
    \top_I.branch[14].l_um_iw[257] ,
    \top_I.branch[14].l_um_iw[256] ,
    \top_I.branch[14].l_um_iw[255] ,
    \top_I.branch[14].l_um_iw[254] ,
    \top_I.branch[14].l_um_iw[253] ,
    \top_I.branch[14].l_um_iw[252] ,
    \top_I.branch[14].l_um_iw[251] ,
    \top_I.branch[14].l_um_iw[250] ,
    \top_I.branch[14].l_um_iw[249] ,
    \top_I.branch[14].l_um_iw[248] ,
    \top_I.branch[14].l_um_iw[247] ,
    \top_I.branch[14].l_um_iw[246] ,
    \top_I.branch[14].l_um_iw[245] ,
    \top_I.branch[14].l_um_iw[244] ,
    \top_I.branch[14].l_um_iw[243] ,
    \top_I.branch[14].l_um_iw[242] ,
    \top_I.branch[14].l_um_iw[241] ,
    \top_I.branch[14].l_um_iw[240] ,
    \top_I.branch[14].l_um_iw[239] ,
    \top_I.branch[14].l_um_iw[238] ,
    \top_I.branch[14].l_um_iw[237] ,
    \top_I.branch[14].l_um_iw[236] ,
    \top_I.branch[14].l_um_iw[235] ,
    \top_I.branch[14].l_um_iw[234] ,
    \top_I.branch[14].l_um_iw[233] ,
    \top_I.branch[14].l_um_iw[232] ,
    \top_I.branch[14].l_um_iw[231] ,
    \top_I.branch[14].l_um_iw[230] ,
    \top_I.branch[14].l_um_iw[229] ,
    \top_I.branch[14].l_um_iw[228] ,
    \top_I.branch[14].l_um_iw[227] ,
    \top_I.branch[14].l_um_iw[226] ,
    \top_I.branch[14].l_um_iw[225] ,
    \top_I.branch[14].l_um_iw[224] ,
    \top_I.branch[14].l_um_iw[223] ,
    \top_I.branch[14].l_um_iw[222] ,
    \top_I.branch[14].l_um_iw[221] ,
    \top_I.branch[14].l_um_iw[220] ,
    \top_I.branch[14].l_um_iw[219] ,
    \top_I.branch[14].l_um_iw[218] ,
    \top_I.branch[14].l_um_iw[217] ,
    \top_I.branch[14].l_um_iw[216] ,
    \top_I.branch[14].l_um_iw[215] ,
    \top_I.branch[14].l_um_iw[214] ,
    \top_I.branch[14].l_um_iw[213] ,
    \top_I.branch[14].l_um_iw[212] ,
    \top_I.branch[14].l_um_iw[211] ,
    \top_I.branch[14].l_um_iw[210] ,
    \top_I.branch[14].l_um_iw[209] ,
    \top_I.branch[14].l_um_iw[208] ,
    \top_I.branch[14].l_um_iw[207] ,
    \top_I.branch[14].l_um_iw[206] ,
    \top_I.branch[14].l_um_iw[205] ,
    \top_I.branch[14].l_um_iw[204] ,
    \top_I.branch[14].l_um_iw[203] ,
    \top_I.branch[14].l_um_iw[202] ,
    \top_I.branch[14].l_um_iw[201] ,
    \top_I.branch[14].l_um_iw[200] ,
    \top_I.branch[14].l_um_iw[199] ,
    \top_I.branch[14].l_um_iw[198] ,
    \top_I.branch[14].l_um_iw[197] ,
    \top_I.branch[14].l_um_iw[196] ,
    \top_I.branch[14].l_um_iw[195] ,
    \top_I.branch[14].l_um_iw[194] ,
    \top_I.branch[14].l_um_iw[193] ,
    \top_I.branch[14].l_um_iw[192] ,
    \top_I.branch[14].l_um_iw[191] ,
    \top_I.branch[14].l_um_iw[190] ,
    \top_I.branch[14].l_um_iw[189] ,
    \top_I.branch[14].l_um_iw[188] ,
    \top_I.branch[14].l_um_iw[187] ,
    \top_I.branch[14].l_um_iw[186] ,
    \top_I.branch[14].l_um_iw[185] ,
    \top_I.branch[14].l_um_iw[184] ,
    \top_I.branch[14].l_um_iw[183] ,
    \top_I.branch[14].l_um_iw[182] ,
    \top_I.branch[14].l_um_iw[181] ,
    \top_I.branch[14].l_um_iw[180] ,
    \top_I.branch[14].l_um_iw[179] ,
    \top_I.branch[14].l_um_iw[178] ,
    \top_I.branch[14].l_um_iw[177] ,
    \top_I.branch[14].l_um_iw[176] ,
    \top_I.branch[14].l_um_iw[175] ,
    \top_I.branch[14].l_um_iw[174] ,
    \top_I.branch[14].l_um_iw[173] ,
    \top_I.branch[14].l_um_iw[172] ,
    \top_I.branch[14].l_um_iw[171] ,
    \top_I.branch[14].l_um_iw[170] ,
    \top_I.branch[14].l_um_iw[169] ,
    \top_I.branch[14].l_um_iw[168] ,
    \top_I.branch[14].l_um_iw[167] ,
    \top_I.branch[14].l_um_iw[166] ,
    \top_I.branch[14].l_um_iw[165] ,
    \top_I.branch[14].l_um_iw[164] ,
    \top_I.branch[14].l_um_iw[163] ,
    \top_I.branch[14].l_um_iw[162] ,
    \top_I.branch[14].l_um_iw[161] ,
    \top_I.branch[14].l_um_iw[160] ,
    \top_I.branch[14].l_um_iw[159] ,
    \top_I.branch[14].l_um_iw[158] ,
    \top_I.branch[14].l_um_iw[157] ,
    \top_I.branch[14].l_um_iw[156] ,
    \top_I.branch[14].l_um_iw[155] ,
    \top_I.branch[14].l_um_iw[154] ,
    \top_I.branch[14].l_um_iw[153] ,
    \top_I.branch[14].l_um_iw[152] ,
    \top_I.branch[14].l_um_iw[151] ,
    \top_I.branch[14].l_um_iw[150] ,
    \top_I.branch[14].l_um_iw[149] ,
    \top_I.branch[14].l_um_iw[148] ,
    \top_I.branch[14].l_um_iw[147] ,
    \top_I.branch[14].l_um_iw[146] ,
    \top_I.branch[14].l_um_iw[145] ,
    \top_I.branch[14].l_um_iw[144] ,
    \top_I.branch[14].l_um_iw[143] ,
    \top_I.branch[14].l_um_iw[142] ,
    \top_I.branch[14].l_um_iw[141] ,
    \top_I.branch[14].l_um_iw[140] ,
    \top_I.branch[14].l_um_iw[139] ,
    \top_I.branch[14].l_um_iw[138] ,
    \top_I.branch[14].l_um_iw[137] ,
    \top_I.branch[14].l_um_iw[136] ,
    \top_I.branch[14].l_um_iw[135] ,
    \top_I.branch[14].l_um_iw[134] ,
    \top_I.branch[14].l_um_iw[133] ,
    \top_I.branch[14].l_um_iw[132] ,
    \top_I.branch[14].l_um_iw[131] ,
    \top_I.branch[14].l_um_iw[130] ,
    \top_I.branch[14].l_um_iw[129] ,
    \top_I.branch[14].l_um_iw[128] ,
    \top_I.branch[14].l_um_iw[127] ,
    \top_I.branch[14].l_um_iw[126] ,
    \top_I.branch[14].l_um_iw[125] ,
    \top_I.branch[14].l_um_iw[124] ,
    \top_I.branch[14].l_um_iw[123] ,
    \top_I.branch[14].l_um_iw[122] ,
    \top_I.branch[14].l_um_iw[121] ,
    \top_I.branch[14].l_um_iw[120] ,
    \top_I.branch[14].l_um_iw[119] ,
    \top_I.branch[14].l_um_iw[118] ,
    \top_I.branch[14].l_um_iw[117] ,
    \top_I.branch[14].l_um_iw[116] ,
    \top_I.branch[14].l_um_iw[115] ,
    \top_I.branch[14].l_um_iw[114] ,
    \top_I.branch[14].l_um_iw[113] ,
    \top_I.branch[14].l_um_iw[112] ,
    \top_I.branch[14].l_um_iw[111] ,
    \top_I.branch[14].l_um_iw[110] ,
    \top_I.branch[14].l_um_iw[109] ,
    \top_I.branch[14].l_um_iw[108] ,
    \top_I.branch[14].l_um_iw[107] ,
    \top_I.branch[14].l_um_iw[106] ,
    \top_I.branch[14].l_um_iw[105] ,
    \top_I.branch[14].l_um_iw[104] ,
    \top_I.branch[14].l_um_iw[103] ,
    \top_I.branch[14].l_um_iw[102] ,
    \top_I.branch[14].l_um_iw[101] ,
    \top_I.branch[14].l_um_iw[100] ,
    \top_I.branch[14].l_um_iw[99] ,
    \top_I.branch[14].l_um_iw[98] ,
    \top_I.branch[14].l_um_iw[97] ,
    \top_I.branch[14].l_um_iw[96] ,
    \top_I.branch[14].l_um_iw[95] ,
    \top_I.branch[14].l_um_iw[94] ,
    \top_I.branch[14].l_um_iw[93] ,
    \top_I.branch[14].l_um_iw[92] ,
    \top_I.branch[14].l_um_iw[91] ,
    \top_I.branch[14].l_um_iw[90] ,
    \top_I.branch[14].l_um_iw[89] ,
    \top_I.branch[14].l_um_iw[88] ,
    \top_I.branch[14].l_um_iw[87] ,
    \top_I.branch[14].l_um_iw[86] ,
    \top_I.branch[14].l_um_iw[85] ,
    \top_I.branch[14].l_um_iw[84] ,
    \top_I.branch[14].l_um_iw[83] ,
    \top_I.branch[14].l_um_iw[82] ,
    \top_I.branch[14].l_um_iw[81] ,
    \top_I.branch[14].l_um_iw[80] ,
    \top_I.branch[14].l_um_iw[79] ,
    \top_I.branch[14].l_um_iw[78] ,
    \top_I.branch[14].l_um_iw[77] ,
    \top_I.branch[14].l_um_iw[76] ,
    \top_I.branch[14].l_um_iw[75] ,
    \top_I.branch[14].l_um_iw[74] ,
    \top_I.branch[14].l_um_iw[73] ,
    \top_I.branch[14].l_um_iw[72] ,
    \top_I.branch[14].l_um_iw[71] ,
    \top_I.branch[14].l_um_iw[70] ,
    \top_I.branch[14].l_um_iw[69] ,
    \top_I.branch[14].l_um_iw[68] ,
    \top_I.branch[14].l_um_iw[67] ,
    \top_I.branch[14].l_um_iw[66] ,
    \top_I.branch[14].l_um_iw[65] ,
    \top_I.branch[14].l_um_iw[64] ,
    \top_I.branch[14].l_um_iw[63] ,
    \top_I.branch[14].l_um_iw[62] ,
    \top_I.branch[14].l_um_iw[61] ,
    \top_I.branch[14].l_um_iw[60] ,
    \top_I.branch[14].l_um_iw[59] ,
    \top_I.branch[14].l_um_iw[58] ,
    \top_I.branch[14].l_um_iw[57] ,
    \top_I.branch[14].l_um_iw[56] ,
    \top_I.branch[14].l_um_iw[55] ,
    \top_I.branch[14].l_um_iw[54] ,
    \top_I.branch[14].l_um_iw[53] ,
    \top_I.branch[14].l_um_iw[52] ,
    \top_I.branch[14].l_um_iw[51] ,
    \top_I.branch[14].l_um_iw[50] ,
    \top_I.branch[14].l_um_iw[49] ,
    \top_I.branch[14].l_um_iw[48] ,
    \top_I.branch[14].l_um_iw[47] ,
    \top_I.branch[14].l_um_iw[46] ,
    \top_I.branch[14].l_um_iw[45] ,
    \top_I.branch[14].l_um_iw[44] ,
    \top_I.branch[14].l_um_iw[43] ,
    \top_I.branch[14].l_um_iw[42] ,
    \top_I.branch[14].l_um_iw[41] ,
    \top_I.branch[14].l_um_iw[40] ,
    \top_I.branch[14].l_um_iw[39] ,
    \top_I.branch[14].l_um_iw[38] ,
    \top_I.branch[14].l_um_iw[37] ,
    \top_I.branch[14].l_um_iw[36] ,
    \top_I.branch[14].l_um_iw[35] ,
    \top_I.branch[14].l_um_iw[34] ,
    \top_I.branch[14].l_um_iw[33] ,
    \top_I.branch[14].l_um_iw[32] ,
    \top_I.branch[14].l_um_iw[31] ,
    \top_I.branch[14].l_um_iw[30] ,
    \top_I.branch[14].l_um_iw[29] ,
    \top_I.branch[14].l_um_iw[28] ,
    \top_I.branch[14].l_um_iw[27] ,
    \top_I.branch[14].l_um_iw[26] ,
    \top_I.branch[14].l_um_iw[25] ,
    \top_I.branch[14].l_um_iw[24] ,
    \top_I.branch[14].l_um_iw[23] ,
    \top_I.branch[14].l_um_iw[22] ,
    \top_I.branch[14].l_um_iw[21] ,
    \top_I.branch[14].l_um_iw[20] ,
    \top_I.branch[14].l_um_iw[19] ,
    \top_I.branch[14].l_um_iw[18] ,
    \top_I.branch[14].l_um_iw[17] ,
    \top_I.branch[14].l_um_iw[16] ,
    \top_I.branch[14].l_um_iw[15] ,
    \top_I.branch[14].l_um_iw[14] ,
    \top_I.branch[14].l_um_iw[13] ,
    \top_I.branch[14].l_um_iw[12] ,
    \top_I.branch[14].l_um_iw[11] ,
    \top_I.branch[14].l_um_iw[10] ,
    \top_I.branch[14].l_um_iw[9] ,
    \top_I.branch[14].l_um_iw[8] ,
    \top_I.branch[14].l_um_iw[7] ,
    \top_I.branch[14].l_um_iw[6] ,
    \top_I.branch[14].l_um_iw[5] ,
    \top_I.branch[14].l_um_iw[4] ,
    \top_I.branch[14].l_um_iw[3] ,
    \top_I.branch[14].l_um_iw[2] ,
    \top_I.branch[14].l_um_iw[1] ,
    \top_I.branch[14].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[1] ,
    \top_I.branch[14].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[15] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[14] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[13] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[12] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[11] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[10] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[9] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[8] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[7] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[6] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[5] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[4] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[3] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].l_um_k_zero[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[14].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] ,
    \top_I.branch[14].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[15].col_um[0].um_top_I.block_15_16.tt_um_I  (.clk(\top_I.branch[15].l_um_iw[18] ),
    .ena(\top_I.branch[15].l_um_ena[1] ),
    .rst_n(\top_I.branch[15].l_um_iw[19] ),
    .ui_in({\top_I.branch[15].l_um_iw[27] ,
    \top_I.branch[15].l_um_iw[26] ,
    \top_I.branch[15].l_um_iw[25] ,
    \top_I.branch[15].l_um_iw[24] ,
    \top_I.branch[15].l_um_iw[23] ,
    \top_I.branch[15].l_um_iw[22] ,
    \top_I.branch[15].l_um_iw[21] ,
    \top_I.branch[15].l_um_iw[20] }),
    .uio_in({\top_I.branch[15].l_um_iw[35] ,
    \top_I.branch[15].l_um_iw[34] ,
    \top_I.branch[15].l_um_iw[33] ,
    \top_I.branch[15].l_um_iw[32] ,
    \top_I.branch[15].l_um_iw[31] ,
    \top_I.branch[15].l_um_iw[30] ,
    \top_I.branch[15].l_um_iw[29] ,
    \top_I.branch[15].l_um_iw[28] }),
    .uio_oe({\top_I.branch[15].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[15].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[15].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[15].mux_I  (.k_one(\top_I.branch[15].l_k_one ),
    .k_zero(\top_I.branch[15].l_k_zero ),
    .addr({\top_I.branch[15].l_k_zero ,
    \top_I.branch[15].l_k_one ,
    \top_I.branch[15].l_k_one ,
    \top_I.branch[15].l_k_one ,
    \top_I.branch[15].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[15].l_um_ena[15] ,
    \top_I.branch[15].l_um_ena[14] ,
    \top_I.branch[15].l_um_ena[13] ,
    \top_I.branch[15].l_um_ena[12] ,
    \top_I.branch[15].l_um_ena[11] ,
    \top_I.branch[15].l_um_ena[10] ,
    \top_I.branch[15].l_um_ena[9] ,
    \top_I.branch[15].l_um_ena[8] ,
    \top_I.branch[15].l_um_ena[7] ,
    \top_I.branch[15].l_um_ena[6] ,
    \top_I.branch[15].l_um_ena[5] ,
    \top_I.branch[15].l_um_ena[4] ,
    \top_I.branch[15].l_um_ena[3] ,
    \top_I.branch[15].l_um_ena[2] ,
    \top_I.branch[15].l_um_ena[1] ,
    \top_I.branch[15].l_um_ena[0] }),
    .um_iw({\top_I.branch[15].l_um_iw[287] ,
    \top_I.branch[15].l_um_iw[286] ,
    \top_I.branch[15].l_um_iw[285] ,
    \top_I.branch[15].l_um_iw[284] ,
    \top_I.branch[15].l_um_iw[283] ,
    \top_I.branch[15].l_um_iw[282] ,
    \top_I.branch[15].l_um_iw[281] ,
    \top_I.branch[15].l_um_iw[280] ,
    \top_I.branch[15].l_um_iw[279] ,
    \top_I.branch[15].l_um_iw[278] ,
    \top_I.branch[15].l_um_iw[277] ,
    \top_I.branch[15].l_um_iw[276] ,
    \top_I.branch[15].l_um_iw[275] ,
    \top_I.branch[15].l_um_iw[274] ,
    \top_I.branch[15].l_um_iw[273] ,
    \top_I.branch[15].l_um_iw[272] ,
    \top_I.branch[15].l_um_iw[271] ,
    \top_I.branch[15].l_um_iw[270] ,
    \top_I.branch[15].l_um_iw[269] ,
    \top_I.branch[15].l_um_iw[268] ,
    \top_I.branch[15].l_um_iw[267] ,
    \top_I.branch[15].l_um_iw[266] ,
    \top_I.branch[15].l_um_iw[265] ,
    \top_I.branch[15].l_um_iw[264] ,
    \top_I.branch[15].l_um_iw[263] ,
    \top_I.branch[15].l_um_iw[262] ,
    \top_I.branch[15].l_um_iw[261] ,
    \top_I.branch[15].l_um_iw[260] ,
    \top_I.branch[15].l_um_iw[259] ,
    \top_I.branch[15].l_um_iw[258] ,
    \top_I.branch[15].l_um_iw[257] ,
    \top_I.branch[15].l_um_iw[256] ,
    \top_I.branch[15].l_um_iw[255] ,
    \top_I.branch[15].l_um_iw[254] ,
    \top_I.branch[15].l_um_iw[253] ,
    \top_I.branch[15].l_um_iw[252] ,
    \top_I.branch[15].l_um_iw[251] ,
    \top_I.branch[15].l_um_iw[250] ,
    \top_I.branch[15].l_um_iw[249] ,
    \top_I.branch[15].l_um_iw[248] ,
    \top_I.branch[15].l_um_iw[247] ,
    \top_I.branch[15].l_um_iw[246] ,
    \top_I.branch[15].l_um_iw[245] ,
    \top_I.branch[15].l_um_iw[244] ,
    \top_I.branch[15].l_um_iw[243] ,
    \top_I.branch[15].l_um_iw[242] ,
    \top_I.branch[15].l_um_iw[241] ,
    \top_I.branch[15].l_um_iw[240] ,
    \top_I.branch[15].l_um_iw[239] ,
    \top_I.branch[15].l_um_iw[238] ,
    \top_I.branch[15].l_um_iw[237] ,
    \top_I.branch[15].l_um_iw[236] ,
    \top_I.branch[15].l_um_iw[235] ,
    \top_I.branch[15].l_um_iw[234] ,
    \top_I.branch[15].l_um_iw[233] ,
    \top_I.branch[15].l_um_iw[232] ,
    \top_I.branch[15].l_um_iw[231] ,
    \top_I.branch[15].l_um_iw[230] ,
    \top_I.branch[15].l_um_iw[229] ,
    \top_I.branch[15].l_um_iw[228] ,
    \top_I.branch[15].l_um_iw[227] ,
    \top_I.branch[15].l_um_iw[226] ,
    \top_I.branch[15].l_um_iw[225] ,
    \top_I.branch[15].l_um_iw[224] ,
    \top_I.branch[15].l_um_iw[223] ,
    \top_I.branch[15].l_um_iw[222] ,
    \top_I.branch[15].l_um_iw[221] ,
    \top_I.branch[15].l_um_iw[220] ,
    \top_I.branch[15].l_um_iw[219] ,
    \top_I.branch[15].l_um_iw[218] ,
    \top_I.branch[15].l_um_iw[217] ,
    \top_I.branch[15].l_um_iw[216] ,
    \top_I.branch[15].l_um_iw[215] ,
    \top_I.branch[15].l_um_iw[214] ,
    \top_I.branch[15].l_um_iw[213] ,
    \top_I.branch[15].l_um_iw[212] ,
    \top_I.branch[15].l_um_iw[211] ,
    \top_I.branch[15].l_um_iw[210] ,
    \top_I.branch[15].l_um_iw[209] ,
    \top_I.branch[15].l_um_iw[208] ,
    \top_I.branch[15].l_um_iw[207] ,
    \top_I.branch[15].l_um_iw[206] ,
    \top_I.branch[15].l_um_iw[205] ,
    \top_I.branch[15].l_um_iw[204] ,
    \top_I.branch[15].l_um_iw[203] ,
    \top_I.branch[15].l_um_iw[202] ,
    \top_I.branch[15].l_um_iw[201] ,
    \top_I.branch[15].l_um_iw[200] ,
    \top_I.branch[15].l_um_iw[199] ,
    \top_I.branch[15].l_um_iw[198] ,
    \top_I.branch[15].l_um_iw[197] ,
    \top_I.branch[15].l_um_iw[196] ,
    \top_I.branch[15].l_um_iw[195] ,
    \top_I.branch[15].l_um_iw[194] ,
    \top_I.branch[15].l_um_iw[193] ,
    \top_I.branch[15].l_um_iw[192] ,
    \top_I.branch[15].l_um_iw[191] ,
    \top_I.branch[15].l_um_iw[190] ,
    \top_I.branch[15].l_um_iw[189] ,
    \top_I.branch[15].l_um_iw[188] ,
    \top_I.branch[15].l_um_iw[187] ,
    \top_I.branch[15].l_um_iw[186] ,
    \top_I.branch[15].l_um_iw[185] ,
    \top_I.branch[15].l_um_iw[184] ,
    \top_I.branch[15].l_um_iw[183] ,
    \top_I.branch[15].l_um_iw[182] ,
    \top_I.branch[15].l_um_iw[181] ,
    \top_I.branch[15].l_um_iw[180] ,
    \top_I.branch[15].l_um_iw[179] ,
    \top_I.branch[15].l_um_iw[178] ,
    \top_I.branch[15].l_um_iw[177] ,
    \top_I.branch[15].l_um_iw[176] ,
    \top_I.branch[15].l_um_iw[175] ,
    \top_I.branch[15].l_um_iw[174] ,
    \top_I.branch[15].l_um_iw[173] ,
    \top_I.branch[15].l_um_iw[172] ,
    \top_I.branch[15].l_um_iw[171] ,
    \top_I.branch[15].l_um_iw[170] ,
    \top_I.branch[15].l_um_iw[169] ,
    \top_I.branch[15].l_um_iw[168] ,
    \top_I.branch[15].l_um_iw[167] ,
    \top_I.branch[15].l_um_iw[166] ,
    \top_I.branch[15].l_um_iw[165] ,
    \top_I.branch[15].l_um_iw[164] ,
    \top_I.branch[15].l_um_iw[163] ,
    \top_I.branch[15].l_um_iw[162] ,
    \top_I.branch[15].l_um_iw[161] ,
    \top_I.branch[15].l_um_iw[160] ,
    \top_I.branch[15].l_um_iw[159] ,
    \top_I.branch[15].l_um_iw[158] ,
    \top_I.branch[15].l_um_iw[157] ,
    \top_I.branch[15].l_um_iw[156] ,
    \top_I.branch[15].l_um_iw[155] ,
    \top_I.branch[15].l_um_iw[154] ,
    \top_I.branch[15].l_um_iw[153] ,
    \top_I.branch[15].l_um_iw[152] ,
    \top_I.branch[15].l_um_iw[151] ,
    \top_I.branch[15].l_um_iw[150] ,
    \top_I.branch[15].l_um_iw[149] ,
    \top_I.branch[15].l_um_iw[148] ,
    \top_I.branch[15].l_um_iw[147] ,
    \top_I.branch[15].l_um_iw[146] ,
    \top_I.branch[15].l_um_iw[145] ,
    \top_I.branch[15].l_um_iw[144] ,
    \top_I.branch[15].l_um_iw[143] ,
    \top_I.branch[15].l_um_iw[142] ,
    \top_I.branch[15].l_um_iw[141] ,
    \top_I.branch[15].l_um_iw[140] ,
    \top_I.branch[15].l_um_iw[139] ,
    \top_I.branch[15].l_um_iw[138] ,
    \top_I.branch[15].l_um_iw[137] ,
    \top_I.branch[15].l_um_iw[136] ,
    \top_I.branch[15].l_um_iw[135] ,
    \top_I.branch[15].l_um_iw[134] ,
    \top_I.branch[15].l_um_iw[133] ,
    \top_I.branch[15].l_um_iw[132] ,
    \top_I.branch[15].l_um_iw[131] ,
    \top_I.branch[15].l_um_iw[130] ,
    \top_I.branch[15].l_um_iw[129] ,
    \top_I.branch[15].l_um_iw[128] ,
    \top_I.branch[15].l_um_iw[127] ,
    \top_I.branch[15].l_um_iw[126] ,
    \top_I.branch[15].l_um_iw[125] ,
    \top_I.branch[15].l_um_iw[124] ,
    \top_I.branch[15].l_um_iw[123] ,
    \top_I.branch[15].l_um_iw[122] ,
    \top_I.branch[15].l_um_iw[121] ,
    \top_I.branch[15].l_um_iw[120] ,
    \top_I.branch[15].l_um_iw[119] ,
    \top_I.branch[15].l_um_iw[118] ,
    \top_I.branch[15].l_um_iw[117] ,
    \top_I.branch[15].l_um_iw[116] ,
    \top_I.branch[15].l_um_iw[115] ,
    \top_I.branch[15].l_um_iw[114] ,
    \top_I.branch[15].l_um_iw[113] ,
    \top_I.branch[15].l_um_iw[112] ,
    \top_I.branch[15].l_um_iw[111] ,
    \top_I.branch[15].l_um_iw[110] ,
    \top_I.branch[15].l_um_iw[109] ,
    \top_I.branch[15].l_um_iw[108] ,
    \top_I.branch[15].l_um_iw[107] ,
    \top_I.branch[15].l_um_iw[106] ,
    \top_I.branch[15].l_um_iw[105] ,
    \top_I.branch[15].l_um_iw[104] ,
    \top_I.branch[15].l_um_iw[103] ,
    \top_I.branch[15].l_um_iw[102] ,
    \top_I.branch[15].l_um_iw[101] ,
    \top_I.branch[15].l_um_iw[100] ,
    \top_I.branch[15].l_um_iw[99] ,
    \top_I.branch[15].l_um_iw[98] ,
    \top_I.branch[15].l_um_iw[97] ,
    \top_I.branch[15].l_um_iw[96] ,
    \top_I.branch[15].l_um_iw[95] ,
    \top_I.branch[15].l_um_iw[94] ,
    \top_I.branch[15].l_um_iw[93] ,
    \top_I.branch[15].l_um_iw[92] ,
    \top_I.branch[15].l_um_iw[91] ,
    \top_I.branch[15].l_um_iw[90] ,
    \top_I.branch[15].l_um_iw[89] ,
    \top_I.branch[15].l_um_iw[88] ,
    \top_I.branch[15].l_um_iw[87] ,
    \top_I.branch[15].l_um_iw[86] ,
    \top_I.branch[15].l_um_iw[85] ,
    \top_I.branch[15].l_um_iw[84] ,
    \top_I.branch[15].l_um_iw[83] ,
    \top_I.branch[15].l_um_iw[82] ,
    \top_I.branch[15].l_um_iw[81] ,
    \top_I.branch[15].l_um_iw[80] ,
    \top_I.branch[15].l_um_iw[79] ,
    \top_I.branch[15].l_um_iw[78] ,
    \top_I.branch[15].l_um_iw[77] ,
    \top_I.branch[15].l_um_iw[76] ,
    \top_I.branch[15].l_um_iw[75] ,
    \top_I.branch[15].l_um_iw[74] ,
    \top_I.branch[15].l_um_iw[73] ,
    \top_I.branch[15].l_um_iw[72] ,
    \top_I.branch[15].l_um_iw[71] ,
    \top_I.branch[15].l_um_iw[70] ,
    \top_I.branch[15].l_um_iw[69] ,
    \top_I.branch[15].l_um_iw[68] ,
    \top_I.branch[15].l_um_iw[67] ,
    \top_I.branch[15].l_um_iw[66] ,
    \top_I.branch[15].l_um_iw[65] ,
    \top_I.branch[15].l_um_iw[64] ,
    \top_I.branch[15].l_um_iw[63] ,
    \top_I.branch[15].l_um_iw[62] ,
    \top_I.branch[15].l_um_iw[61] ,
    \top_I.branch[15].l_um_iw[60] ,
    \top_I.branch[15].l_um_iw[59] ,
    \top_I.branch[15].l_um_iw[58] ,
    \top_I.branch[15].l_um_iw[57] ,
    \top_I.branch[15].l_um_iw[56] ,
    \top_I.branch[15].l_um_iw[55] ,
    \top_I.branch[15].l_um_iw[54] ,
    \top_I.branch[15].l_um_iw[53] ,
    \top_I.branch[15].l_um_iw[52] ,
    \top_I.branch[15].l_um_iw[51] ,
    \top_I.branch[15].l_um_iw[50] ,
    \top_I.branch[15].l_um_iw[49] ,
    \top_I.branch[15].l_um_iw[48] ,
    \top_I.branch[15].l_um_iw[47] ,
    \top_I.branch[15].l_um_iw[46] ,
    \top_I.branch[15].l_um_iw[45] ,
    \top_I.branch[15].l_um_iw[44] ,
    \top_I.branch[15].l_um_iw[43] ,
    \top_I.branch[15].l_um_iw[42] ,
    \top_I.branch[15].l_um_iw[41] ,
    \top_I.branch[15].l_um_iw[40] ,
    \top_I.branch[15].l_um_iw[39] ,
    \top_I.branch[15].l_um_iw[38] ,
    \top_I.branch[15].l_um_iw[37] ,
    \top_I.branch[15].l_um_iw[36] ,
    \top_I.branch[15].l_um_iw[35] ,
    \top_I.branch[15].l_um_iw[34] ,
    \top_I.branch[15].l_um_iw[33] ,
    \top_I.branch[15].l_um_iw[32] ,
    \top_I.branch[15].l_um_iw[31] ,
    \top_I.branch[15].l_um_iw[30] ,
    \top_I.branch[15].l_um_iw[29] ,
    \top_I.branch[15].l_um_iw[28] ,
    \top_I.branch[15].l_um_iw[27] ,
    \top_I.branch[15].l_um_iw[26] ,
    \top_I.branch[15].l_um_iw[25] ,
    \top_I.branch[15].l_um_iw[24] ,
    \top_I.branch[15].l_um_iw[23] ,
    \top_I.branch[15].l_um_iw[22] ,
    \top_I.branch[15].l_um_iw[21] ,
    \top_I.branch[15].l_um_iw[20] ,
    \top_I.branch[15].l_um_iw[19] ,
    \top_I.branch[15].l_um_iw[18] ,
    \top_I.branch[15].l_um_iw[17] ,
    \top_I.branch[15].l_um_iw[16] ,
    \top_I.branch[15].l_um_iw[15] ,
    \top_I.branch[15].l_um_iw[14] ,
    \top_I.branch[15].l_um_iw[13] ,
    \top_I.branch[15].l_um_iw[12] ,
    \top_I.branch[15].l_um_iw[11] ,
    \top_I.branch[15].l_um_iw[10] ,
    \top_I.branch[15].l_um_iw[9] ,
    \top_I.branch[15].l_um_iw[8] ,
    \top_I.branch[15].l_um_iw[7] ,
    \top_I.branch[15].l_um_iw[6] ,
    \top_I.branch[15].l_um_iw[5] ,
    \top_I.branch[15].l_um_iw[4] ,
    \top_I.branch[15].l_um_iw[3] ,
    \top_I.branch[15].l_um_iw[2] ,
    \top_I.branch[15].l_um_iw[1] ,
    \top_I.branch[15].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[1] ,
    \top_I.branch[15].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[15] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[14] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[13] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[12] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[11] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[10] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[9] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[8] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[7] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[6] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[5] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[4] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[3] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].l_um_k_zero[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[15].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] ,
    \top_I.branch[15].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[16].col_um[0].um_bot_I.block_16_0.tt_um_I  (.clk(\top_I.branch[16].l_um_iw[0] ),
    .ena(\top_I.branch[16].l_um_ena[0] ),
    .rst_n(\top_I.branch[16].l_um_iw[1] ),
    .ui_in({\top_I.branch[16].l_um_iw[9] ,
    \top_I.branch[16].l_um_iw[8] ,
    \top_I.branch[16].l_um_iw[7] ,
    \top_I.branch[16].l_um_iw[6] ,
    \top_I.branch[16].l_um_iw[5] ,
    \top_I.branch[16].l_um_iw[4] ,
    \top_I.branch[16].l_um_iw[3] ,
    \top_I.branch[16].l_um_iw[2] }),
    .uio_in({\top_I.branch[16].l_um_iw[17] ,
    \top_I.branch[16].l_um_iw[16] ,
    \top_I.branch[16].l_um_iw[15] ,
    \top_I.branch[16].l_um_iw[14] ,
    \top_I.branch[16].l_um_iw[13] ,
    \top_I.branch[16].l_um_iw[12] ,
    \top_I.branch[16].l_um_iw[11] ,
    \top_I.branch[16].l_um_iw[10] }),
    .uio_oe({\top_I.branch[16].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[16].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[16].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[16].mux_I  (.k_one(\top_I.branch[16].l_k_one ),
    .k_zero(\top_I.branch[16].l_k_zero ),
    .addr({\top_I.branch[16].l_k_one ,
    \top_I.branch[16].l_k_zero ,
    \top_I.branch[16].l_k_zero ,
    \top_I.branch[16].l_k_zero ,
    \top_I.branch[16].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[16].l_um_ena[15] ,
    \top_I.branch[16].l_um_ena[14] ,
    \top_I.branch[16].l_um_ena[13] ,
    \top_I.branch[16].l_um_ena[12] ,
    \top_I.branch[16].l_um_ena[11] ,
    \top_I.branch[16].l_um_ena[10] ,
    \top_I.branch[16].l_um_ena[9] ,
    \top_I.branch[16].l_um_ena[8] ,
    \top_I.branch[16].l_um_ena[7] ,
    \top_I.branch[16].l_um_ena[6] ,
    \top_I.branch[16].l_um_ena[5] ,
    \top_I.branch[16].l_um_ena[4] ,
    \top_I.branch[16].l_um_ena[3] ,
    \top_I.branch[16].l_um_ena[2] ,
    \top_I.branch[16].l_um_ena[1] ,
    \top_I.branch[16].l_um_ena[0] }),
    .um_iw({\top_I.branch[16].l_um_iw[287] ,
    \top_I.branch[16].l_um_iw[286] ,
    \top_I.branch[16].l_um_iw[285] ,
    \top_I.branch[16].l_um_iw[284] ,
    \top_I.branch[16].l_um_iw[283] ,
    \top_I.branch[16].l_um_iw[282] ,
    \top_I.branch[16].l_um_iw[281] ,
    \top_I.branch[16].l_um_iw[280] ,
    \top_I.branch[16].l_um_iw[279] ,
    \top_I.branch[16].l_um_iw[278] ,
    \top_I.branch[16].l_um_iw[277] ,
    \top_I.branch[16].l_um_iw[276] ,
    \top_I.branch[16].l_um_iw[275] ,
    \top_I.branch[16].l_um_iw[274] ,
    \top_I.branch[16].l_um_iw[273] ,
    \top_I.branch[16].l_um_iw[272] ,
    \top_I.branch[16].l_um_iw[271] ,
    \top_I.branch[16].l_um_iw[270] ,
    \top_I.branch[16].l_um_iw[269] ,
    \top_I.branch[16].l_um_iw[268] ,
    \top_I.branch[16].l_um_iw[267] ,
    \top_I.branch[16].l_um_iw[266] ,
    \top_I.branch[16].l_um_iw[265] ,
    \top_I.branch[16].l_um_iw[264] ,
    \top_I.branch[16].l_um_iw[263] ,
    \top_I.branch[16].l_um_iw[262] ,
    \top_I.branch[16].l_um_iw[261] ,
    \top_I.branch[16].l_um_iw[260] ,
    \top_I.branch[16].l_um_iw[259] ,
    \top_I.branch[16].l_um_iw[258] ,
    \top_I.branch[16].l_um_iw[257] ,
    \top_I.branch[16].l_um_iw[256] ,
    \top_I.branch[16].l_um_iw[255] ,
    \top_I.branch[16].l_um_iw[254] ,
    \top_I.branch[16].l_um_iw[253] ,
    \top_I.branch[16].l_um_iw[252] ,
    \top_I.branch[16].l_um_iw[251] ,
    \top_I.branch[16].l_um_iw[250] ,
    \top_I.branch[16].l_um_iw[249] ,
    \top_I.branch[16].l_um_iw[248] ,
    \top_I.branch[16].l_um_iw[247] ,
    \top_I.branch[16].l_um_iw[246] ,
    \top_I.branch[16].l_um_iw[245] ,
    \top_I.branch[16].l_um_iw[244] ,
    \top_I.branch[16].l_um_iw[243] ,
    \top_I.branch[16].l_um_iw[242] ,
    \top_I.branch[16].l_um_iw[241] ,
    \top_I.branch[16].l_um_iw[240] ,
    \top_I.branch[16].l_um_iw[239] ,
    \top_I.branch[16].l_um_iw[238] ,
    \top_I.branch[16].l_um_iw[237] ,
    \top_I.branch[16].l_um_iw[236] ,
    \top_I.branch[16].l_um_iw[235] ,
    \top_I.branch[16].l_um_iw[234] ,
    \top_I.branch[16].l_um_iw[233] ,
    \top_I.branch[16].l_um_iw[232] ,
    \top_I.branch[16].l_um_iw[231] ,
    \top_I.branch[16].l_um_iw[230] ,
    \top_I.branch[16].l_um_iw[229] ,
    \top_I.branch[16].l_um_iw[228] ,
    \top_I.branch[16].l_um_iw[227] ,
    \top_I.branch[16].l_um_iw[226] ,
    \top_I.branch[16].l_um_iw[225] ,
    \top_I.branch[16].l_um_iw[224] ,
    \top_I.branch[16].l_um_iw[223] ,
    \top_I.branch[16].l_um_iw[222] ,
    \top_I.branch[16].l_um_iw[221] ,
    \top_I.branch[16].l_um_iw[220] ,
    \top_I.branch[16].l_um_iw[219] ,
    \top_I.branch[16].l_um_iw[218] ,
    \top_I.branch[16].l_um_iw[217] ,
    \top_I.branch[16].l_um_iw[216] ,
    \top_I.branch[16].l_um_iw[215] ,
    \top_I.branch[16].l_um_iw[214] ,
    \top_I.branch[16].l_um_iw[213] ,
    \top_I.branch[16].l_um_iw[212] ,
    \top_I.branch[16].l_um_iw[211] ,
    \top_I.branch[16].l_um_iw[210] ,
    \top_I.branch[16].l_um_iw[209] ,
    \top_I.branch[16].l_um_iw[208] ,
    \top_I.branch[16].l_um_iw[207] ,
    \top_I.branch[16].l_um_iw[206] ,
    \top_I.branch[16].l_um_iw[205] ,
    \top_I.branch[16].l_um_iw[204] ,
    \top_I.branch[16].l_um_iw[203] ,
    \top_I.branch[16].l_um_iw[202] ,
    \top_I.branch[16].l_um_iw[201] ,
    \top_I.branch[16].l_um_iw[200] ,
    \top_I.branch[16].l_um_iw[199] ,
    \top_I.branch[16].l_um_iw[198] ,
    \top_I.branch[16].l_um_iw[197] ,
    \top_I.branch[16].l_um_iw[196] ,
    \top_I.branch[16].l_um_iw[195] ,
    \top_I.branch[16].l_um_iw[194] ,
    \top_I.branch[16].l_um_iw[193] ,
    \top_I.branch[16].l_um_iw[192] ,
    \top_I.branch[16].l_um_iw[191] ,
    \top_I.branch[16].l_um_iw[190] ,
    \top_I.branch[16].l_um_iw[189] ,
    \top_I.branch[16].l_um_iw[188] ,
    \top_I.branch[16].l_um_iw[187] ,
    \top_I.branch[16].l_um_iw[186] ,
    \top_I.branch[16].l_um_iw[185] ,
    \top_I.branch[16].l_um_iw[184] ,
    \top_I.branch[16].l_um_iw[183] ,
    \top_I.branch[16].l_um_iw[182] ,
    \top_I.branch[16].l_um_iw[181] ,
    \top_I.branch[16].l_um_iw[180] ,
    \top_I.branch[16].l_um_iw[179] ,
    \top_I.branch[16].l_um_iw[178] ,
    \top_I.branch[16].l_um_iw[177] ,
    \top_I.branch[16].l_um_iw[176] ,
    \top_I.branch[16].l_um_iw[175] ,
    \top_I.branch[16].l_um_iw[174] ,
    \top_I.branch[16].l_um_iw[173] ,
    \top_I.branch[16].l_um_iw[172] ,
    \top_I.branch[16].l_um_iw[171] ,
    \top_I.branch[16].l_um_iw[170] ,
    \top_I.branch[16].l_um_iw[169] ,
    \top_I.branch[16].l_um_iw[168] ,
    \top_I.branch[16].l_um_iw[167] ,
    \top_I.branch[16].l_um_iw[166] ,
    \top_I.branch[16].l_um_iw[165] ,
    \top_I.branch[16].l_um_iw[164] ,
    \top_I.branch[16].l_um_iw[163] ,
    \top_I.branch[16].l_um_iw[162] ,
    \top_I.branch[16].l_um_iw[161] ,
    \top_I.branch[16].l_um_iw[160] ,
    \top_I.branch[16].l_um_iw[159] ,
    \top_I.branch[16].l_um_iw[158] ,
    \top_I.branch[16].l_um_iw[157] ,
    \top_I.branch[16].l_um_iw[156] ,
    \top_I.branch[16].l_um_iw[155] ,
    \top_I.branch[16].l_um_iw[154] ,
    \top_I.branch[16].l_um_iw[153] ,
    \top_I.branch[16].l_um_iw[152] ,
    \top_I.branch[16].l_um_iw[151] ,
    \top_I.branch[16].l_um_iw[150] ,
    \top_I.branch[16].l_um_iw[149] ,
    \top_I.branch[16].l_um_iw[148] ,
    \top_I.branch[16].l_um_iw[147] ,
    \top_I.branch[16].l_um_iw[146] ,
    \top_I.branch[16].l_um_iw[145] ,
    \top_I.branch[16].l_um_iw[144] ,
    \top_I.branch[16].l_um_iw[143] ,
    \top_I.branch[16].l_um_iw[142] ,
    \top_I.branch[16].l_um_iw[141] ,
    \top_I.branch[16].l_um_iw[140] ,
    \top_I.branch[16].l_um_iw[139] ,
    \top_I.branch[16].l_um_iw[138] ,
    \top_I.branch[16].l_um_iw[137] ,
    \top_I.branch[16].l_um_iw[136] ,
    \top_I.branch[16].l_um_iw[135] ,
    \top_I.branch[16].l_um_iw[134] ,
    \top_I.branch[16].l_um_iw[133] ,
    \top_I.branch[16].l_um_iw[132] ,
    \top_I.branch[16].l_um_iw[131] ,
    \top_I.branch[16].l_um_iw[130] ,
    \top_I.branch[16].l_um_iw[129] ,
    \top_I.branch[16].l_um_iw[128] ,
    \top_I.branch[16].l_um_iw[127] ,
    \top_I.branch[16].l_um_iw[126] ,
    \top_I.branch[16].l_um_iw[125] ,
    \top_I.branch[16].l_um_iw[124] ,
    \top_I.branch[16].l_um_iw[123] ,
    \top_I.branch[16].l_um_iw[122] ,
    \top_I.branch[16].l_um_iw[121] ,
    \top_I.branch[16].l_um_iw[120] ,
    \top_I.branch[16].l_um_iw[119] ,
    \top_I.branch[16].l_um_iw[118] ,
    \top_I.branch[16].l_um_iw[117] ,
    \top_I.branch[16].l_um_iw[116] ,
    \top_I.branch[16].l_um_iw[115] ,
    \top_I.branch[16].l_um_iw[114] ,
    \top_I.branch[16].l_um_iw[113] ,
    \top_I.branch[16].l_um_iw[112] ,
    \top_I.branch[16].l_um_iw[111] ,
    \top_I.branch[16].l_um_iw[110] ,
    \top_I.branch[16].l_um_iw[109] ,
    \top_I.branch[16].l_um_iw[108] ,
    \top_I.branch[16].l_um_iw[107] ,
    \top_I.branch[16].l_um_iw[106] ,
    \top_I.branch[16].l_um_iw[105] ,
    \top_I.branch[16].l_um_iw[104] ,
    \top_I.branch[16].l_um_iw[103] ,
    \top_I.branch[16].l_um_iw[102] ,
    \top_I.branch[16].l_um_iw[101] ,
    \top_I.branch[16].l_um_iw[100] ,
    \top_I.branch[16].l_um_iw[99] ,
    \top_I.branch[16].l_um_iw[98] ,
    \top_I.branch[16].l_um_iw[97] ,
    \top_I.branch[16].l_um_iw[96] ,
    \top_I.branch[16].l_um_iw[95] ,
    \top_I.branch[16].l_um_iw[94] ,
    \top_I.branch[16].l_um_iw[93] ,
    \top_I.branch[16].l_um_iw[92] ,
    \top_I.branch[16].l_um_iw[91] ,
    \top_I.branch[16].l_um_iw[90] ,
    \top_I.branch[16].l_um_iw[89] ,
    \top_I.branch[16].l_um_iw[88] ,
    \top_I.branch[16].l_um_iw[87] ,
    \top_I.branch[16].l_um_iw[86] ,
    \top_I.branch[16].l_um_iw[85] ,
    \top_I.branch[16].l_um_iw[84] ,
    \top_I.branch[16].l_um_iw[83] ,
    \top_I.branch[16].l_um_iw[82] ,
    \top_I.branch[16].l_um_iw[81] ,
    \top_I.branch[16].l_um_iw[80] ,
    \top_I.branch[16].l_um_iw[79] ,
    \top_I.branch[16].l_um_iw[78] ,
    \top_I.branch[16].l_um_iw[77] ,
    \top_I.branch[16].l_um_iw[76] ,
    \top_I.branch[16].l_um_iw[75] ,
    \top_I.branch[16].l_um_iw[74] ,
    \top_I.branch[16].l_um_iw[73] ,
    \top_I.branch[16].l_um_iw[72] ,
    \top_I.branch[16].l_um_iw[71] ,
    \top_I.branch[16].l_um_iw[70] ,
    \top_I.branch[16].l_um_iw[69] ,
    \top_I.branch[16].l_um_iw[68] ,
    \top_I.branch[16].l_um_iw[67] ,
    \top_I.branch[16].l_um_iw[66] ,
    \top_I.branch[16].l_um_iw[65] ,
    \top_I.branch[16].l_um_iw[64] ,
    \top_I.branch[16].l_um_iw[63] ,
    \top_I.branch[16].l_um_iw[62] ,
    \top_I.branch[16].l_um_iw[61] ,
    \top_I.branch[16].l_um_iw[60] ,
    \top_I.branch[16].l_um_iw[59] ,
    \top_I.branch[16].l_um_iw[58] ,
    \top_I.branch[16].l_um_iw[57] ,
    \top_I.branch[16].l_um_iw[56] ,
    \top_I.branch[16].l_um_iw[55] ,
    \top_I.branch[16].l_um_iw[54] ,
    \top_I.branch[16].l_um_iw[53] ,
    \top_I.branch[16].l_um_iw[52] ,
    \top_I.branch[16].l_um_iw[51] ,
    \top_I.branch[16].l_um_iw[50] ,
    \top_I.branch[16].l_um_iw[49] ,
    \top_I.branch[16].l_um_iw[48] ,
    \top_I.branch[16].l_um_iw[47] ,
    \top_I.branch[16].l_um_iw[46] ,
    \top_I.branch[16].l_um_iw[45] ,
    \top_I.branch[16].l_um_iw[44] ,
    \top_I.branch[16].l_um_iw[43] ,
    \top_I.branch[16].l_um_iw[42] ,
    \top_I.branch[16].l_um_iw[41] ,
    \top_I.branch[16].l_um_iw[40] ,
    \top_I.branch[16].l_um_iw[39] ,
    \top_I.branch[16].l_um_iw[38] ,
    \top_I.branch[16].l_um_iw[37] ,
    \top_I.branch[16].l_um_iw[36] ,
    \top_I.branch[16].l_um_iw[35] ,
    \top_I.branch[16].l_um_iw[34] ,
    \top_I.branch[16].l_um_iw[33] ,
    \top_I.branch[16].l_um_iw[32] ,
    \top_I.branch[16].l_um_iw[31] ,
    \top_I.branch[16].l_um_iw[30] ,
    \top_I.branch[16].l_um_iw[29] ,
    \top_I.branch[16].l_um_iw[28] ,
    \top_I.branch[16].l_um_iw[27] ,
    \top_I.branch[16].l_um_iw[26] ,
    \top_I.branch[16].l_um_iw[25] ,
    \top_I.branch[16].l_um_iw[24] ,
    \top_I.branch[16].l_um_iw[23] ,
    \top_I.branch[16].l_um_iw[22] ,
    \top_I.branch[16].l_um_iw[21] ,
    \top_I.branch[16].l_um_iw[20] ,
    \top_I.branch[16].l_um_iw[19] ,
    \top_I.branch[16].l_um_iw[18] ,
    \top_I.branch[16].l_um_iw[17] ,
    \top_I.branch[16].l_um_iw[16] ,
    \top_I.branch[16].l_um_iw[15] ,
    \top_I.branch[16].l_um_iw[14] ,
    \top_I.branch[16].l_um_iw[13] ,
    \top_I.branch[16].l_um_iw[12] ,
    \top_I.branch[16].l_um_iw[11] ,
    \top_I.branch[16].l_um_iw[10] ,
    \top_I.branch[16].l_um_iw[9] ,
    \top_I.branch[16].l_um_iw[8] ,
    \top_I.branch[16].l_um_iw[7] ,
    \top_I.branch[16].l_um_iw[6] ,
    \top_I.branch[16].l_um_iw[5] ,
    \top_I.branch[16].l_um_iw[4] ,
    \top_I.branch[16].l_um_iw[3] ,
    \top_I.branch[16].l_um_iw[2] ,
    \top_I.branch[16].l_um_iw[1] ,
    \top_I.branch[16].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[15] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[14] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[13] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[12] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[11] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[10] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[9] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[8] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[7] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[6] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[5] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[4] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[3] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[2] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].l_um_k_zero[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[16].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[17].col_um[0].um_bot_I.block_16_16.tt_um_I  (.clk(\top_I.branch[17].l_um_iw[0] ),
    .ena(\top_I.branch[17].l_um_ena[0] ),
    .rst_n(\top_I.branch[17].l_um_iw[1] ),
    .ui_in({\top_I.branch[17].l_um_iw[9] ,
    \top_I.branch[17].l_um_iw[8] ,
    \top_I.branch[17].l_um_iw[7] ,
    \top_I.branch[17].l_um_iw[6] ,
    \top_I.branch[17].l_um_iw[5] ,
    \top_I.branch[17].l_um_iw[4] ,
    \top_I.branch[17].l_um_iw[3] ,
    \top_I.branch[17].l_um_iw[2] }),
    .uio_in({\top_I.branch[17].l_um_iw[17] ,
    \top_I.branch[17].l_um_iw[16] ,
    \top_I.branch[17].l_um_iw[15] ,
    \top_I.branch[17].l_um_iw[14] ,
    \top_I.branch[17].l_um_iw[13] ,
    \top_I.branch[17].l_um_iw[12] ,
    \top_I.branch[17].l_um_iw[11] ,
    \top_I.branch[17].l_um_iw[10] }),
    .uio_oe({\top_I.branch[17].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[17].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[17].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[17].mux_I  (.k_one(\top_I.branch[17].l_k_one ),
    .k_zero(\top_I.branch[17].l_k_zero ),
    .addr({\top_I.branch[17].l_k_one ,
    \top_I.branch[17].l_k_zero ,
    \top_I.branch[17].l_k_zero ,
    \top_I.branch[17].l_k_zero ,
    \top_I.branch[17].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[17].l_um_ena[15] ,
    \top_I.branch[17].l_um_ena[14] ,
    \top_I.branch[17].l_um_ena[13] ,
    \top_I.branch[17].l_um_ena[12] ,
    \top_I.branch[17].l_um_ena[11] ,
    \top_I.branch[17].l_um_ena[10] ,
    \top_I.branch[17].l_um_ena[9] ,
    \top_I.branch[17].l_um_ena[8] ,
    \top_I.branch[17].l_um_ena[7] ,
    \top_I.branch[17].l_um_ena[6] ,
    \top_I.branch[17].l_um_ena[5] ,
    \top_I.branch[17].l_um_ena[4] ,
    \top_I.branch[17].l_um_ena[3] ,
    \top_I.branch[17].l_um_ena[2] ,
    \top_I.branch[17].l_um_ena[1] ,
    \top_I.branch[17].l_um_ena[0] }),
    .um_iw({\top_I.branch[17].l_um_iw[287] ,
    \top_I.branch[17].l_um_iw[286] ,
    \top_I.branch[17].l_um_iw[285] ,
    \top_I.branch[17].l_um_iw[284] ,
    \top_I.branch[17].l_um_iw[283] ,
    \top_I.branch[17].l_um_iw[282] ,
    \top_I.branch[17].l_um_iw[281] ,
    \top_I.branch[17].l_um_iw[280] ,
    \top_I.branch[17].l_um_iw[279] ,
    \top_I.branch[17].l_um_iw[278] ,
    \top_I.branch[17].l_um_iw[277] ,
    \top_I.branch[17].l_um_iw[276] ,
    \top_I.branch[17].l_um_iw[275] ,
    \top_I.branch[17].l_um_iw[274] ,
    \top_I.branch[17].l_um_iw[273] ,
    \top_I.branch[17].l_um_iw[272] ,
    \top_I.branch[17].l_um_iw[271] ,
    \top_I.branch[17].l_um_iw[270] ,
    \top_I.branch[17].l_um_iw[269] ,
    \top_I.branch[17].l_um_iw[268] ,
    \top_I.branch[17].l_um_iw[267] ,
    \top_I.branch[17].l_um_iw[266] ,
    \top_I.branch[17].l_um_iw[265] ,
    \top_I.branch[17].l_um_iw[264] ,
    \top_I.branch[17].l_um_iw[263] ,
    \top_I.branch[17].l_um_iw[262] ,
    \top_I.branch[17].l_um_iw[261] ,
    \top_I.branch[17].l_um_iw[260] ,
    \top_I.branch[17].l_um_iw[259] ,
    \top_I.branch[17].l_um_iw[258] ,
    \top_I.branch[17].l_um_iw[257] ,
    \top_I.branch[17].l_um_iw[256] ,
    \top_I.branch[17].l_um_iw[255] ,
    \top_I.branch[17].l_um_iw[254] ,
    \top_I.branch[17].l_um_iw[253] ,
    \top_I.branch[17].l_um_iw[252] ,
    \top_I.branch[17].l_um_iw[251] ,
    \top_I.branch[17].l_um_iw[250] ,
    \top_I.branch[17].l_um_iw[249] ,
    \top_I.branch[17].l_um_iw[248] ,
    \top_I.branch[17].l_um_iw[247] ,
    \top_I.branch[17].l_um_iw[246] ,
    \top_I.branch[17].l_um_iw[245] ,
    \top_I.branch[17].l_um_iw[244] ,
    \top_I.branch[17].l_um_iw[243] ,
    \top_I.branch[17].l_um_iw[242] ,
    \top_I.branch[17].l_um_iw[241] ,
    \top_I.branch[17].l_um_iw[240] ,
    \top_I.branch[17].l_um_iw[239] ,
    \top_I.branch[17].l_um_iw[238] ,
    \top_I.branch[17].l_um_iw[237] ,
    \top_I.branch[17].l_um_iw[236] ,
    \top_I.branch[17].l_um_iw[235] ,
    \top_I.branch[17].l_um_iw[234] ,
    \top_I.branch[17].l_um_iw[233] ,
    \top_I.branch[17].l_um_iw[232] ,
    \top_I.branch[17].l_um_iw[231] ,
    \top_I.branch[17].l_um_iw[230] ,
    \top_I.branch[17].l_um_iw[229] ,
    \top_I.branch[17].l_um_iw[228] ,
    \top_I.branch[17].l_um_iw[227] ,
    \top_I.branch[17].l_um_iw[226] ,
    \top_I.branch[17].l_um_iw[225] ,
    \top_I.branch[17].l_um_iw[224] ,
    \top_I.branch[17].l_um_iw[223] ,
    \top_I.branch[17].l_um_iw[222] ,
    \top_I.branch[17].l_um_iw[221] ,
    \top_I.branch[17].l_um_iw[220] ,
    \top_I.branch[17].l_um_iw[219] ,
    \top_I.branch[17].l_um_iw[218] ,
    \top_I.branch[17].l_um_iw[217] ,
    \top_I.branch[17].l_um_iw[216] ,
    \top_I.branch[17].l_um_iw[215] ,
    \top_I.branch[17].l_um_iw[214] ,
    \top_I.branch[17].l_um_iw[213] ,
    \top_I.branch[17].l_um_iw[212] ,
    \top_I.branch[17].l_um_iw[211] ,
    \top_I.branch[17].l_um_iw[210] ,
    \top_I.branch[17].l_um_iw[209] ,
    \top_I.branch[17].l_um_iw[208] ,
    \top_I.branch[17].l_um_iw[207] ,
    \top_I.branch[17].l_um_iw[206] ,
    \top_I.branch[17].l_um_iw[205] ,
    \top_I.branch[17].l_um_iw[204] ,
    \top_I.branch[17].l_um_iw[203] ,
    \top_I.branch[17].l_um_iw[202] ,
    \top_I.branch[17].l_um_iw[201] ,
    \top_I.branch[17].l_um_iw[200] ,
    \top_I.branch[17].l_um_iw[199] ,
    \top_I.branch[17].l_um_iw[198] ,
    \top_I.branch[17].l_um_iw[197] ,
    \top_I.branch[17].l_um_iw[196] ,
    \top_I.branch[17].l_um_iw[195] ,
    \top_I.branch[17].l_um_iw[194] ,
    \top_I.branch[17].l_um_iw[193] ,
    \top_I.branch[17].l_um_iw[192] ,
    \top_I.branch[17].l_um_iw[191] ,
    \top_I.branch[17].l_um_iw[190] ,
    \top_I.branch[17].l_um_iw[189] ,
    \top_I.branch[17].l_um_iw[188] ,
    \top_I.branch[17].l_um_iw[187] ,
    \top_I.branch[17].l_um_iw[186] ,
    \top_I.branch[17].l_um_iw[185] ,
    \top_I.branch[17].l_um_iw[184] ,
    \top_I.branch[17].l_um_iw[183] ,
    \top_I.branch[17].l_um_iw[182] ,
    \top_I.branch[17].l_um_iw[181] ,
    \top_I.branch[17].l_um_iw[180] ,
    \top_I.branch[17].l_um_iw[179] ,
    \top_I.branch[17].l_um_iw[178] ,
    \top_I.branch[17].l_um_iw[177] ,
    \top_I.branch[17].l_um_iw[176] ,
    \top_I.branch[17].l_um_iw[175] ,
    \top_I.branch[17].l_um_iw[174] ,
    \top_I.branch[17].l_um_iw[173] ,
    \top_I.branch[17].l_um_iw[172] ,
    \top_I.branch[17].l_um_iw[171] ,
    \top_I.branch[17].l_um_iw[170] ,
    \top_I.branch[17].l_um_iw[169] ,
    \top_I.branch[17].l_um_iw[168] ,
    \top_I.branch[17].l_um_iw[167] ,
    \top_I.branch[17].l_um_iw[166] ,
    \top_I.branch[17].l_um_iw[165] ,
    \top_I.branch[17].l_um_iw[164] ,
    \top_I.branch[17].l_um_iw[163] ,
    \top_I.branch[17].l_um_iw[162] ,
    \top_I.branch[17].l_um_iw[161] ,
    \top_I.branch[17].l_um_iw[160] ,
    \top_I.branch[17].l_um_iw[159] ,
    \top_I.branch[17].l_um_iw[158] ,
    \top_I.branch[17].l_um_iw[157] ,
    \top_I.branch[17].l_um_iw[156] ,
    \top_I.branch[17].l_um_iw[155] ,
    \top_I.branch[17].l_um_iw[154] ,
    \top_I.branch[17].l_um_iw[153] ,
    \top_I.branch[17].l_um_iw[152] ,
    \top_I.branch[17].l_um_iw[151] ,
    \top_I.branch[17].l_um_iw[150] ,
    \top_I.branch[17].l_um_iw[149] ,
    \top_I.branch[17].l_um_iw[148] ,
    \top_I.branch[17].l_um_iw[147] ,
    \top_I.branch[17].l_um_iw[146] ,
    \top_I.branch[17].l_um_iw[145] ,
    \top_I.branch[17].l_um_iw[144] ,
    \top_I.branch[17].l_um_iw[143] ,
    \top_I.branch[17].l_um_iw[142] ,
    \top_I.branch[17].l_um_iw[141] ,
    \top_I.branch[17].l_um_iw[140] ,
    \top_I.branch[17].l_um_iw[139] ,
    \top_I.branch[17].l_um_iw[138] ,
    \top_I.branch[17].l_um_iw[137] ,
    \top_I.branch[17].l_um_iw[136] ,
    \top_I.branch[17].l_um_iw[135] ,
    \top_I.branch[17].l_um_iw[134] ,
    \top_I.branch[17].l_um_iw[133] ,
    \top_I.branch[17].l_um_iw[132] ,
    \top_I.branch[17].l_um_iw[131] ,
    \top_I.branch[17].l_um_iw[130] ,
    \top_I.branch[17].l_um_iw[129] ,
    \top_I.branch[17].l_um_iw[128] ,
    \top_I.branch[17].l_um_iw[127] ,
    \top_I.branch[17].l_um_iw[126] ,
    \top_I.branch[17].l_um_iw[125] ,
    \top_I.branch[17].l_um_iw[124] ,
    \top_I.branch[17].l_um_iw[123] ,
    \top_I.branch[17].l_um_iw[122] ,
    \top_I.branch[17].l_um_iw[121] ,
    \top_I.branch[17].l_um_iw[120] ,
    \top_I.branch[17].l_um_iw[119] ,
    \top_I.branch[17].l_um_iw[118] ,
    \top_I.branch[17].l_um_iw[117] ,
    \top_I.branch[17].l_um_iw[116] ,
    \top_I.branch[17].l_um_iw[115] ,
    \top_I.branch[17].l_um_iw[114] ,
    \top_I.branch[17].l_um_iw[113] ,
    \top_I.branch[17].l_um_iw[112] ,
    \top_I.branch[17].l_um_iw[111] ,
    \top_I.branch[17].l_um_iw[110] ,
    \top_I.branch[17].l_um_iw[109] ,
    \top_I.branch[17].l_um_iw[108] ,
    \top_I.branch[17].l_um_iw[107] ,
    \top_I.branch[17].l_um_iw[106] ,
    \top_I.branch[17].l_um_iw[105] ,
    \top_I.branch[17].l_um_iw[104] ,
    \top_I.branch[17].l_um_iw[103] ,
    \top_I.branch[17].l_um_iw[102] ,
    \top_I.branch[17].l_um_iw[101] ,
    \top_I.branch[17].l_um_iw[100] ,
    \top_I.branch[17].l_um_iw[99] ,
    \top_I.branch[17].l_um_iw[98] ,
    \top_I.branch[17].l_um_iw[97] ,
    \top_I.branch[17].l_um_iw[96] ,
    \top_I.branch[17].l_um_iw[95] ,
    \top_I.branch[17].l_um_iw[94] ,
    \top_I.branch[17].l_um_iw[93] ,
    \top_I.branch[17].l_um_iw[92] ,
    \top_I.branch[17].l_um_iw[91] ,
    \top_I.branch[17].l_um_iw[90] ,
    \top_I.branch[17].l_um_iw[89] ,
    \top_I.branch[17].l_um_iw[88] ,
    \top_I.branch[17].l_um_iw[87] ,
    \top_I.branch[17].l_um_iw[86] ,
    \top_I.branch[17].l_um_iw[85] ,
    \top_I.branch[17].l_um_iw[84] ,
    \top_I.branch[17].l_um_iw[83] ,
    \top_I.branch[17].l_um_iw[82] ,
    \top_I.branch[17].l_um_iw[81] ,
    \top_I.branch[17].l_um_iw[80] ,
    \top_I.branch[17].l_um_iw[79] ,
    \top_I.branch[17].l_um_iw[78] ,
    \top_I.branch[17].l_um_iw[77] ,
    \top_I.branch[17].l_um_iw[76] ,
    \top_I.branch[17].l_um_iw[75] ,
    \top_I.branch[17].l_um_iw[74] ,
    \top_I.branch[17].l_um_iw[73] ,
    \top_I.branch[17].l_um_iw[72] ,
    \top_I.branch[17].l_um_iw[71] ,
    \top_I.branch[17].l_um_iw[70] ,
    \top_I.branch[17].l_um_iw[69] ,
    \top_I.branch[17].l_um_iw[68] ,
    \top_I.branch[17].l_um_iw[67] ,
    \top_I.branch[17].l_um_iw[66] ,
    \top_I.branch[17].l_um_iw[65] ,
    \top_I.branch[17].l_um_iw[64] ,
    \top_I.branch[17].l_um_iw[63] ,
    \top_I.branch[17].l_um_iw[62] ,
    \top_I.branch[17].l_um_iw[61] ,
    \top_I.branch[17].l_um_iw[60] ,
    \top_I.branch[17].l_um_iw[59] ,
    \top_I.branch[17].l_um_iw[58] ,
    \top_I.branch[17].l_um_iw[57] ,
    \top_I.branch[17].l_um_iw[56] ,
    \top_I.branch[17].l_um_iw[55] ,
    \top_I.branch[17].l_um_iw[54] ,
    \top_I.branch[17].l_um_iw[53] ,
    \top_I.branch[17].l_um_iw[52] ,
    \top_I.branch[17].l_um_iw[51] ,
    \top_I.branch[17].l_um_iw[50] ,
    \top_I.branch[17].l_um_iw[49] ,
    \top_I.branch[17].l_um_iw[48] ,
    \top_I.branch[17].l_um_iw[47] ,
    \top_I.branch[17].l_um_iw[46] ,
    \top_I.branch[17].l_um_iw[45] ,
    \top_I.branch[17].l_um_iw[44] ,
    \top_I.branch[17].l_um_iw[43] ,
    \top_I.branch[17].l_um_iw[42] ,
    \top_I.branch[17].l_um_iw[41] ,
    \top_I.branch[17].l_um_iw[40] ,
    \top_I.branch[17].l_um_iw[39] ,
    \top_I.branch[17].l_um_iw[38] ,
    \top_I.branch[17].l_um_iw[37] ,
    \top_I.branch[17].l_um_iw[36] ,
    \top_I.branch[17].l_um_iw[35] ,
    \top_I.branch[17].l_um_iw[34] ,
    \top_I.branch[17].l_um_iw[33] ,
    \top_I.branch[17].l_um_iw[32] ,
    \top_I.branch[17].l_um_iw[31] ,
    \top_I.branch[17].l_um_iw[30] ,
    \top_I.branch[17].l_um_iw[29] ,
    \top_I.branch[17].l_um_iw[28] ,
    \top_I.branch[17].l_um_iw[27] ,
    \top_I.branch[17].l_um_iw[26] ,
    \top_I.branch[17].l_um_iw[25] ,
    \top_I.branch[17].l_um_iw[24] ,
    \top_I.branch[17].l_um_iw[23] ,
    \top_I.branch[17].l_um_iw[22] ,
    \top_I.branch[17].l_um_iw[21] ,
    \top_I.branch[17].l_um_iw[20] ,
    \top_I.branch[17].l_um_iw[19] ,
    \top_I.branch[17].l_um_iw[18] ,
    \top_I.branch[17].l_um_iw[17] ,
    \top_I.branch[17].l_um_iw[16] ,
    \top_I.branch[17].l_um_iw[15] ,
    \top_I.branch[17].l_um_iw[14] ,
    \top_I.branch[17].l_um_iw[13] ,
    \top_I.branch[17].l_um_iw[12] ,
    \top_I.branch[17].l_um_iw[11] ,
    \top_I.branch[17].l_um_iw[10] ,
    \top_I.branch[17].l_um_iw[9] ,
    \top_I.branch[17].l_um_iw[8] ,
    \top_I.branch[17].l_um_iw[7] ,
    \top_I.branch[17].l_um_iw[6] ,
    \top_I.branch[17].l_um_iw[5] ,
    \top_I.branch[17].l_um_iw[4] ,
    \top_I.branch[17].l_um_iw[3] ,
    \top_I.branch[17].l_um_iw[2] ,
    \top_I.branch[17].l_um_iw[1] ,
    \top_I.branch[17].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[15] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[14] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[13] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[12] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[11] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[10] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[9] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[8] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[7] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[6] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[5] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[4] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[3] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[2] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].l_um_k_zero[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[17].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[18].col_um[0].um_top_I.block_19_0.tt_um_I  (.clk(\top_I.branch[18].l_um_iw[18] ),
    .ena(\top_I.branch[18].l_um_ena[1] ),
    .rst_n(\top_I.branch[18].l_um_iw[19] ),
    .ui_in({\top_I.branch[18].l_um_iw[27] ,
    \top_I.branch[18].l_um_iw[26] ,
    \top_I.branch[18].l_um_iw[25] ,
    \top_I.branch[18].l_um_iw[24] ,
    \top_I.branch[18].l_um_iw[23] ,
    \top_I.branch[18].l_um_iw[22] ,
    \top_I.branch[18].l_um_iw[21] ,
    \top_I.branch[18].l_um_iw[20] }),
    .uio_in({\top_I.branch[18].l_um_iw[35] ,
    \top_I.branch[18].l_um_iw[34] ,
    \top_I.branch[18].l_um_iw[33] ,
    \top_I.branch[18].l_um_iw[32] ,
    \top_I.branch[18].l_um_iw[31] ,
    \top_I.branch[18].l_um_iw[30] ,
    \top_I.branch[18].l_um_iw[29] ,
    \top_I.branch[18].l_um_iw[28] }),
    .uio_oe({\top_I.branch[18].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[18].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[18].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[18].mux_I  (.k_one(\top_I.branch[18].l_k_one ),
    .k_zero(\top_I.branch[18].l_k_zero ),
    .addr({\top_I.branch[18].l_k_one ,
    \top_I.branch[18].l_k_zero ,
    \top_I.branch[18].l_k_zero ,
    \top_I.branch[18].l_k_one ,
    \top_I.branch[18].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[18].l_um_ena[15] ,
    \top_I.branch[18].l_um_ena[14] ,
    \top_I.branch[18].l_um_ena[13] ,
    \top_I.branch[18].l_um_ena[12] ,
    \top_I.branch[18].l_um_ena[11] ,
    \top_I.branch[18].l_um_ena[10] ,
    \top_I.branch[18].l_um_ena[9] ,
    \top_I.branch[18].l_um_ena[8] ,
    \top_I.branch[18].l_um_ena[7] ,
    \top_I.branch[18].l_um_ena[6] ,
    \top_I.branch[18].l_um_ena[5] ,
    \top_I.branch[18].l_um_ena[4] ,
    \top_I.branch[18].l_um_ena[3] ,
    \top_I.branch[18].l_um_ena[2] ,
    \top_I.branch[18].l_um_ena[1] ,
    \top_I.branch[18].l_um_ena[0] }),
    .um_iw({\top_I.branch[18].l_um_iw[287] ,
    \top_I.branch[18].l_um_iw[286] ,
    \top_I.branch[18].l_um_iw[285] ,
    \top_I.branch[18].l_um_iw[284] ,
    \top_I.branch[18].l_um_iw[283] ,
    \top_I.branch[18].l_um_iw[282] ,
    \top_I.branch[18].l_um_iw[281] ,
    \top_I.branch[18].l_um_iw[280] ,
    \top_I.branch[18].l_um_iw[279] ,
    \top_I.branch[18].l_um_iw[278] ,
    \top_I.branch[18].l_um_iw[277] ,
    \top_I.branch[18].l_um_iw[276] ,
    \top_I.branch[18].l_um_iw[275] ,
    \top_I.branch[18].l_um_iw[274] ,
    \top_I.branch[18].l_um_iw[273] ,
    \top_I.branch[18].l_um_iw[272] ,
    \top_I.branch[18].l_um_iw[271] ,
    \top_I.branch[18].l_um_iw[270] ,
    \top_I.branch[18].l_um_iw[269] ,
    \top_I.branch[18].l_um_iw[268] ,
    \top_I.branch[18].l_um_iw[267] ,
    \top_I.branch[18].l_um_iw[266] ,
    \top_I.branch[18].l_um_iw[265] ,
    \top_I.branch[18].l_um_iw[264] ,
    \top_I.branch[18].l_um_iw[263] ,
    \top_I.branch[18].l_um_iw[262] ,
    \top_I.branch[18].l_um_iw[261] ,
    \top_I.branch[18].l_um_iw[260] ,
    \top_I.branch[18].l_um_iw[259] ,
    \top_I.branch[18].l_um_iw[258] ,
    \top_I.branch[18].l_um_iw[257] ,
    \top_I.branch[18].l_um_iw[256] ,
    \top_I.branch[18].l_um_iw[255] ,
    \top_I.branch[18].l_um_iw[254] ,
    \top_I.branch[18].l_um_iw[253] ,
    \top_I.branch[18].l_um_iw[252] ,
    \top_I.branch[18].l_um_iw[251] ,
    \top_I.branch[18].l_um_iw[250] ,
    \top_I.branch[18].l_um_iw[249] ,
    \top_I.branch[18].l_um_iw[248] ,
    \top_I.branch[18].l_um_iw[247] ,
    \top_I.branch[18].l_um_iw[246] ,
    \top_I.branch[18].l_um_iw[245] ,
    \top_I.branch[18].l_um_iw[244] ,
    \top_I.branch[18].l_um_iw[243] ,
    \top_I.branch[18].l_um_iw[242] ,
    \top_I.branch[18].l_um_iw[241] ,
    \top_I.branch[18].l_um_iw[240] ,
    \top_I.branch[18].l_um_iw[239] ,
    \top_I.branch[18].l_um_iw[238] ,
    \top_I.branch[18].l_um_iw[237] ,
    \top_I.branch[18].l_um_iw[236] ,
    \top_I.branch[18].l_um_iw[235] ,
    \top_I.branch[18].l_um_iw[234] ,
    \top_I.branch[18].l_um_iw[233] ,
    \top_I.branch[18].l_um_iw[232] ,
    \top_I.branch[18].l_um_iw[231] ,
    \top_I.branch[18].l_um_iw[230] ,
    \top_I.branch[18].l_um_iw[229] ,
    \top_I.branch[18].l_um_iw[228] ,
    \top_I.branch[18].l_um_iw[227] ,
    \top_I.branch[18].l_um_iw[226] ,
    \top_I.branch[18].l_um_iw[225] ,
    \top_I.branch[18].l_um_iw[224] ,
    \top_I.branch[18].l_um_iw[223] ,
    \top_I.branch[18].l_um_iw[222] ,
    \top_I.branch[18].l_um_iw[221] ,
    \top_I.branch[18].l_um_iw[220] ,
    \top_I.branch[18].l_um_iw[219] ,
    \top_I.branch[18].l_um_iw[218] ,
    \top_I.branch[18].l_um_iw[217] ,
    \top_I.branch[18].l_um_iw[216] ,
    \top_I.branch[18].l_um_iw[215] ,
    \top_I.branch[18].l_um_iw[214] ,
    \top_I.branch[18].l_um_iw[213] ,
    \top_I.branch[18].l_um_iw[212] ,
    \top_I.branch[18].l_um_iw[211] ,
    \top_I.branch[18].l_um_iw[210] ,
    \top_I.branch[18].l_um_iw[209] ,
    \top_I.branch[18].l_um_iw[208] ,
    \top_I.branch[18].l_um_iw[207] ,
    \top_I.branch[18].l_um_iw[206] ,
    \top_I.branch[18].l_um_iw[205] ,
    \top_I.branch[18].l_um_iw[204] ,
    \top_I.branch[18].l_um_iw[203] ,
    \top_I.branch[18].l_um_iw[202] ,
    \top_I.branch[18].l_um_iw[201] ,
    \top_I.branch[18].l_um_iw[200] ,
    \top_I.branch[18].l_um_iw[199] ,
    \top_I.branch[18].l_um_iw[198] ,
    \top_I.branch[18].l_um_iw[197] ,
    \top_I.branch[18].l_um_iw[196] ,
    \top_I.branch[18].l_um_iw[195] ,
    \top_I.branch[18].l_um_iw[194] ,
    \top_I.branch[18].l_um_iw[193] ,
    \top_I.branch[18].l_um_iw[192] ,
    \top_I.branch[18].l_um_iw[191] ,
    \top_I.branch[18].l_um_iw[190] ,
    \top_I.branch[18].l_um_iw[189] ,
    \top_I.branch[18].l_um_iw[188] ,
    \top_I.branch[18].l_um_iw[187] ,
    \top_I.branch[18].l_um_iw[186] ,
    \top_I.branch[18].l_um_iw[185] ,
    \top_I.branch[18].l_um_iw[184] ,
    \top_I.branch[18].l_um_iw[183] ,
    \top_I.branch[18].l_um_iw[182] ,
    \top_I.branch[18].l_um_iw[181] ,
    \top_I.branch[18].l_um_iw[180] ,
    \top_I.branch[18].l_um_iw[179] ,
    \top_I.branch[18].l_um_iw[178] ,
    \top_I.branch[18].l_um_iw[177] ,
    \top_I.branch[18].l_um_iw[176] ,
    \top_I.branch[18].l_um_iw[175] ,
    \top_I.branch[18].l_um_iw[174] ,
    \top_I.branch[18].l_um_iw[173] ,
    \top_I.branch[18].l_um_iw[172] ,
    \top_I.branch[18].l_um_iw[171] ,
    \top_I.branch[18].l_um_iw[170] ,
    \top_I.branch[18].l_um_iw[169] ,
    \top_I.branch[18].l_um_iw[168] ,
    \top_I.branch[18].l_um_iw[167] ,
    \top_I.branch[18].l_um_iw[166] ,
    \top_I.branch[18].l_um_iw[165] ,
    \top_I.branch[18].l_um_iw[164] ,
    \top_I.branch[18].l_um_iw[163] ,
    \top_I.branch[18].l_um_iw[162] ,
    \top_I.branch[18].l_um_iw[161] ,
    \top_I.branch[18].l_um_iw[160] ,
    \top_I.branch[18].l_um_iw[159] ,
    \top_I.branch[18].l_um_iw[158] ,
    \top_I.branch[18].l_um_iw[157] ,
    \top_I.branch[18].l_um_iw[156] ,
    \top_I.branch[18].l_um_iw[155] ,
    \top_I.branch[18].l_um_iw[154] ,
    \top_I.branch[18].l_um_iw[153] ,
    \top_I.branch[18].l_um_iw[152] ,
    \top_I.branch[18].l_um_iw[151] ,
    \top_I.branch[18].l_um_iw[150] ,
    \top_I.branch[18].l_um_iw[149] ,
    \top_I.branch[18].l_um_iw[148] ,
    \top_I.branch[18].l_um_iw[147] ,
    \top_I.branch[18].l_um_iw[146] ,
    \top_I.branch[18].l_um_iw[145] ,
    \top_I.branch[18].l_um_iw[144] ,
    \top_I.branch[18].l_um_iw[143] ,
    \top_I.branch[18].l_um_iw[142] ,
    \top_I.branch[18].l_um_iw[141] ,
    \top_I.branch[18].l_um_iw[140] ,
    \top_I.branch[18].l_um_iw[139] ,
    \top_I.branch[18].l_um_iw[138] ,
    \top_I.branch[18].l_um_iw[137] ,
    \top_I.branch[18].l_um_iw[136] ,
    \top_I.branch[18].l_um_iw[135] ,
    \top_I.branch[18].l_um_iw[134] ,
    \top_I.branch[18].l_um_iw[133] ,
    \top_I.branch[18].l_um_iw[132] ,
    \top_I.branch[18].l_um_iw[131] ,
    \top_I.branch[18].l_um_iw[130] ,
    \top_I.branch[18].l_um_iw[129] ,
    \top_I.branch[18].l_um_iw[128] ,
    \top_I.branch[18].l_um_iw[127] ,
    \top_I.branch[18].l_um_iw[126] ,
    \top_I.branch[18].l_um_iw[125] ,
    \top_I.branch[18].l_um_iw[124] ,
    \top_I.branch[18].l_um_iw[123] ,
    \top_I.branch[18].l_um_iw[122] ,
    \top_I.branch[18].l_um_iw[121] ,
    \top_I.branch[18].l_um_iw[120] ,
    \top_I.branch[18].l_um_iw[119] ,
    \top_I.branch[18].l_um_iw[118] ,
    \top_I.branch[18].l_um_iw[117] ,
    \top_I.branch[18].l_um_iw[116] ,
    \top_I.branch[18].l_um_iw[115] ,
    \top_I.branch[18].l_um_iw[114] ,
    \top_I.branch[18].l_um_iw[113] ,
    \top_I.branch[18].l_um_iw[112] ,
    \top_I.branch[18].l_um_iw[111] ,
    \top_I.branch[18].l_um_iw[110] ,
    \top_I.branch[18].l_um_iw[109] ,
    \top_I.branch[18].l_um_iw[108] ,
    \top_I.branch[18].l_um_iw[107] ,
    \top_I.branch[18].l_um_iw[106] ,
    \top_I.branch[18].l_um_iw[105] ,
    \top_I.branch[18].l_um_iw[104] ,
    \top_I.branch[18].l_um_iw[103] ,
    \top_I.branch[18].l_um_iw[102] ,
    \top_I.branch[18].l_um_iw[101] ,
    \top_I.branch[18].l_um_iw[100] ,
    \top_I.branch[18].l_um_iw[99] ,
    \top_I.branch[18].l_um_iw[98] ,
    \top_I.branch[18].l_um_iw[97] ,
    \top_I.branch[18].l_um_iw[96] ,
    \top_I.branch[18].l_um_iw[95] ,
    \top_I.branch[18].l_um_iw[94] ,
    \top_I.branch[18].l_um_iw[93] ,
    \top_I.branch[18].l_um_iw[92] ,
    \top_I.branch[18].l_um_iw[91] ,
    \top_I.branch[18].l_um_iw[90] ,
    \top_I.branch[18].l_um_iw[89] ,
    \top_I.branch[18].l_um_iw[88] ,
    \top_I.branch[18].l_um_iw[87] ,
    \top_I.branch[18].l_um_iw[86] ,
    \top_I.branch[18].l_um_iw[85] ,
    \top_I.branch[18].l_um_iw[84] ,
    \top_I.branch[18].l_um_iw[83] ,
    \top_I.branch[18].l_um_iw[82] ,
    \top_I.branch[18].l_um_iw[81] ,
    \top_I.branch[18].l_um_iw[80] ,
    \top_I.branch[18].l_um_iw[79] ,
    \top_I.branch[18].l_um_iw[78] ,
    \top_I.branch[18].l_um_iw[77] ,
    \top_I.branch[18].l_um_iw[76] ,
    \top_I.branch[18].l_um_iw[75] ,
    \top_I.branch[18].l_um_iw[74] ,
    \top_I.branch[18].l_um_iw[73] ,
    \top_I.branch[18].l_um_iw[72] ,
    \top_I.branch[18].l_um_iw[71] ,
    \top_I.branch[18].l_um_iw[70] ,
    \top_I.branch[18].l_um_iw[69] ,
    \top_I.branch[18].l_um_iw[68] ,
    \top_I.branch[18].l_um_iw[67] ,
    \top_I.branch[18].l_um_iw[66] ,
    \top_I.branch[18].l_um_iw[65] ,
    \top_I.branch[18].l_um_iw[64] ,
    \top_I.branch[18].l_um_iw[63] ,
    \top_I.branch[18].l_um_iw[62] ,
    \top_I.branch[18].l_um_iw[61] ,
    \top_I.branch[18].l_um_iw[60] ,
    \top_I.branch[18].l_um_iw[59] ,
    \top_I.branch[18].l_um_iw[58] ,
    \top_I.branch[18].l_um_iw[57] ,
    \top_I.branch[18].l_um_iw[56] ,
    \top_I.branch[18].l_um_iw[55] ,
    \top_I.branch[18].l_um_iw[54] ,
    \top_I.branch[18].l_um_iw[53] ,
    \top_I.branch[18].l_um_iw[52] ,
    \top_I.branch[18].l_um_iw[51] ,
    \top_I.branch[18].l_um_iw[50] ,
    \top_I.branch[18].l_um_iw[49] ,
    \top_I.branch[18].l_um_iw[48] ,
    \top_I.branch[18].l_um_iw[47] ,
    \top_I.branch[18].l_um_iw[46] ,
    \top_I.branch[18].l_um_iw[45] ,
    \top_I.branch[18].l_um_iw[44] ,
    \top_I.branch[18].l_um_iw[43] ,
    \top_I.branch[18].l_um_iw[42] ,
    \top_I.branch[18].l_um_iw[41] ,
    \top_I.branch[18].l_um_iw[40] ,
    \top_I.branch[18].l_um_iw[39] ,
    \top_I.branch[18].l_um_iw[38] ,
    \top_I.branch[18].l_um_iw[37] ,
    \top_I.branch[18].l_um_iw[36] ,
    \top_I.branch[18].l_um_iw[35] ,
    \top_I.branch[18].l_um_iw[34] ,
    \top_I.branch[18].l_um_iw[33] ,
    \top_I.branch[18].l_um_iw[32] ,
    \top_I.branch[18].l_um_iw[31] ,
    \top_I.branch[18].l_um_iw[30] ,
    \top_I.branch[18].l_um_iw[29] ,
    \top_I.branch[18].l_um_iw[28] ,
    \top_I.branch[18].l_um_iw[27] ,
    \top_I.branch[18].l_um_iw[26] ,
    \top_I.branch[18].l_um_iw[25] ,
    \top_I.branch[18].l_um_iw[24] ,
    \top_I.branch[18].l_um_iw[23] ,
    \top_I.branch[18].l_um_iw[22] ,
    \top_I.branch[18].l_um_iw[21] ,
    \top_I.branch[18].l_um_iw[20] ,
    \top_I.branch[18].l_um_iw[19] ,
    \top_I.branch[18].l_um_iw[18] ,
    \top_I.branch[18].l_um_iw[17] ,
    \top_I.branch[18].l_um_iw[16] ,
    \top_I.branch[18].l_um_iw[15] ,
    \top_I.branch[18].l_um_iw[14] ,
    \top_I.branch[18].l_um_iw[13] ,
    \top_I.branch[18].l_um_iw[12] ,
    \top_I.branch[18].l_um_iw[11] ,
    \top_I.branch[18].l_um_iw[10] ,
    \top_I.branch[18].l_um_iw[9] ,
    \top_I.branch[18].l_um_iw[8] ,
    \top_I.branch[18].l_um_iw[7] ,
    \top_I.branch[18].l_um_iw[6] ,
    \top_I.branch[18].l_um_iw[5] ,
    \top_I.branch[18].l_um_iw[4] ,
    \top_I.branch[18].l_um_iw[3] ,
    \top_I.branch[18].l_um_iw[2] ,
    \top_I.branch[18].l_um_iw[1] ,
    \top_I.branch[18].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[1] ,
    \top_I.branch[18].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[15] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[14] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[13] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[12] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[11] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[10] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[9] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[8] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[7] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[6] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[5] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[4] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[3] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].l_um_k_zero[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[18].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] ,
    \top_I.branch[18].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[19].col_um[0].um_top_I.block_19_16.tt_um_I  (.clk(\top_I.branch[19].l_um_iw[18] ),
    .ena(\top_I.branch[19].l_um_ena[1] ),
    .rst_n(\top_I.branch[19].l_um_iw[19] ),
    .ui_in({\top_I.branch[19].l_um_iw[27] ,
    \top_I.branch[19].l_um_iw[26] ,
    \top_I.branch[19].l_um_iw[25] ,
    \top_I.branch[19].l_um_iw[24] ,
    \top_I.branch[19].l_um_iw[23] ,
    \top_I.branch[19].l_um_iw[22] ,
    \top_I.branch[19].l_um_iw[21] ,
    \top_I.branch[19].l_um_iw[20] }),
    .uio_in({\top_I.branch[19].l_um_iw[35] ,
    \top_I.branch[19].l_um_iw[34] ,
    \top_I.branch[19].l_um_iw[33] ,
    \top_I.branch[19].l_um_iw[32] ,
    \top_I.branch[19].l_um_iw[31] ,
    \top_I.branch[19].l_um_iw[30] ,
    \top_I.branch[19].l_um_iw[29] ,
    \top_I.branch[19].l_um_iw[28] }),
    .uio_oe({\top_I.branch[19].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[19].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[19].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[19].mux_I  (.k_one(\top_I.branch[19].l_k_one ),
    .k_zero(\top_I.branch[19].l_k_zero ),
    .addr({\top_I.branch[19].l_k_one ,
    \top_I.branch[19].l_k_zero ,
    \top_I.branch[19].l_k_zero ,
    \top_I.branch[19].l_k_one ,
    \top_I.branch[19].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[19].l_um_ena[15] ,
    \top_I.branch[19].l_um_ena[14] ,
    \top_I.branch[19].l_um_ena[13] ,
    \top_I.branch[19].l_um_ena[12] ,
    \top_I.branch[19].l_um_ena[11] ,
    \top_I.branch[19].l_um_ena[10] ,
    \top_I.branch[19].l_um_ena[9] ,
    \top_I.branch[19].l_um_ena[8] ,
    \top_I.branch[19].l_um_ena[7] ,
    \top_I.branch[19].l_um_ena[6] ,
    \top_I.branch[19].l_um_ena[5] ,
    \top_I.branch[19].l_um_ena[4] ,
    \top_I.branch[19].l_um_ena[3] ,
    \top_I.branch[19].l_um_ena[2] ,
    \top_I.branch[19].l_um_ena[1] ,
    \top_I.branch[19].l_um_ena[0] }),
    .um_iw({\top_I.branch[19].l_um_iw[287] ,
    \top_I.branch[19].l_um_iw[286] ,
    \top_I.branch[19].l_um_iw[285] ,
    \top_I.branch[19].l_um_iw[284] ,
    \top_I.branch[19].l_um_iw[283] ,
    \top_I.branch[19].l_um_iw[282] ,
    \top_I.branch[19].l_um_iw[281] ,
    \top_I.branch[19].l_um_iw[280] ,
    \top_I.branch[19].l_um_iw[279] ,
    \top_I.branch[19].l_um_iw[278] ,
    \top_I.branch[19].l_um_iw[277] ,
    \top_I.branch[19].l_um_iw[276] ,
    \top_I.branch[19].l_um_iw[275] ,
    \top_I.branch[19].l_um_iw[274] ,
    \top_I.branch[19].l_um_iw[273] ,
    \top_I.branch[19].l_um_iw[272] ,
    \top_I.branch[19].l_um_iw[271] ,
    \top_I.branch[19].l_um_iw[270] ,
    \top_I.branch[19].l_um_iw[269] ,
    \top_I.branch[19].l_um_iw[268] ,
    \top_I.branch[19].l_um_iw[267] ,
    \top_I.branch[19].l_um_iw[266] ,
    \top_I.branch[19].l_um_iw[265] ,
    \top_I.branch[19].l_um_iw[264] ,
    \top_I.branch[19].l_um_iw[263] ,
    \top_I.branch[19].l_um_iw[262] ,
    \top_I.branch[19].l_um_iw[261] ,
    \top_I.branch[19].l_um_iw[260] ,
    \top_I.branch[19].l_um_iw[259] ,
    \top_I.branch[19].l_um_iw[258] ,
    \top_I.branch[19].l_um_iw[257] ,
    \top_I.branch[19].l_um_iw[256] ,
    \top_I.branch[19].l_um_iw[255] ,
    \top_I.branch[19].l_um_iw[254] ,
    \top_I.branch[19].l_um_iw[253] ,
    \top_I.branch[19].l_um_iw[252] ,
    \top_I.branch[19].l_um_iw[251] ,
    \top_I.branch[19].l_um_iw[250] ,
    \top_I.branch[19].l_um_iw[249] ,
    \top_I.branch[19].l_um_iw[248] ,
    \top_I.branch[19].l_um_iw[247] ,
    \top_I.branch[19].l_um_iw[246] ,
    \top_I.branch[19].l_um_iw[245] ,
    \top_I.branch[19].l_um_iw[244] ,
    \top_I.branch[19].l_um_iw[243] ,
    \top_I.branch[19].l_um_iw[242] ,
    \top_I.branch[19].l_um_iw[241] ,
    \top_I.branch[19].l_um_iw[240] ,
    \top_I.branch[19].l_um_iw[239] ,
    \top_I.branch[19].l_um_iw[238] ,
    \top_I.branch[19].l_um_iw[237] ,
    \top_I.branch[19].l_um_iw[236] ,
    \top_I.branch[19].l_um_iw[235] ,
    \top_I.branch[19].l_um_iw[234] ,
    \top_I.branch[19].l_um_iw[233] ,
    \top_I.branch[19].l_um_iw[232] ,
    \top_I.branch[19].l_um_iw[231] ,
    \top_I.branch[19].l_um_iw[230] ,
    \top_I.branch[19].l_um_iw[229] ,
    \top_I.branch[19].l_um_iw[228] ,
    \top_I.branch[19].l_um_iw[227] ,
    \top_I.branch[19].l_um_iw[226] ,
    \top_I.branch[19].l_um_iw[225] ,
    \top_I.branch[19].l_um_iw[224] ,
    \top_I.branch[19].l_um_iw[223] ,
    \top_I.branch[19].l_um_iw[222] ,
    \top_I.branch[19].l_um_iw[221] ,
    \top_I.branch[19].l_um_iw[220] ,
    \top_I.branch[19].l_um_iw[219] ,
    \top_I.branch[19].l_um_iw[218] ,
    \top_I.branch[19].l_um_iw[217] ,
    \top_I.branch[19].l_um_iw[216] ,
    \top_I.branch[19].l_um_iw[215] ,
    \top_I.branch[19].l_um_iw[214] ,
    \top_I.branch[19].l_um_iw[213] ,
    \top_I.branch[19].l_um_iw[212] ,
    \top_I.branch[19].l_um_iw[211] ,
    \top_I.branch[19].l_um_iw[210] ,
    \top_I.branch[19].l_um_iw[209] ,
    \top_I.branch[19].l_um_iw[208] ,
    \top_I.branch[19].l_um_iw[207] ,
    \top_I.branch[19].l_um_iw[206] ,
    \top_I.branch[19].l_um_iw[205] ,
    \top_I.branch[19].l_um_iw[204] ,
    \top_I.branch[19].l_um_iw[203] ,
    \top_I.branch[19].l_um_iw[202] ,
    \top_I.branch[19].l_um_iw[201] ,
    \top_I.branch[19].l_um_iw[200] ,
    \top_I.branch[19].l_um_iw[199] ,
    \top_I.branch[19].l_um_iw[198] ,
    \top_I.branch[19].l_um_iw[197] ,
    \top_I.branch[19].l_um_iw[196] ,
    \top_I.branch[19].l_um_iw[195] ,
    \top_I.branch[19].l_um_iw[194] ,
    \top_I.branch[19].l_um_iw[193] ,
    \top_I.branch[19].l_um_iw[192] ,
    \top_I.branch[19].l_um_iw[191] ,
    \top_I.branch[19].l_um_iw[190] ,
    \top_I.branch[19].l_um_iw[189] ,
    \top_I.branch[19].l_um_iw[188] ,
    \top_I.branch[19].l_um_iw[187] ,
    \top_I.branch[19].l_um_iw[186] ,
    \top_I.branch[19].l_um_iw[185] ,
    \top_I.branch[19].l_um_iw[184] ,
    \top_I.branch[19].l_um_iw[183] ,
    \top_I.branch[19].l_um_iw[182] ,
    \top_I.branch[19].l_um_iw[181] ,
    \top_I.branch[19].l_um_iw[180] ,
    \top_I.branch[19].l_um_iw[179] ,
    \top_I.branch[19].l_um_iw[178] ,
    \top_I.branch[19].l_um_iw[177] ,
    \top_I.branch[19].l_um_iw[176] ,
    \top_I.branch[19].l_um_iw[175] ,
    \top_I.branch[19].l_um_iw[174] ,
    \top_I.branch[19].l_um_iw[173] ,
    \top_I.branch[19].l_um_iw[172] ,
    \top_I.branch[19].l_um_iw[171] ,
    \top_I.branch[19].l_um_iw[170] ,
    \top_I.branch[19].l_um_iw[169] ,
    \top_I.branch[19].l_um_iw[168] ,
    \top_I.branch[19].l_um_iw[167] ,
    \top_I.branch[19].l_um_iw[166] ,
    \top_I.branch[19].l_um_iw[165] ,
    \top_I.branch[19].l_um_iw[164] ,
    \top_I.branch[19].l_um_iw[163] ,
    \top_I.branch[19].l_um_iw[162] ,
    \top_I.branch[19].l_um_iw[161] ,
    \top_I.branch[19].l_um_iw[160] ,
    \top_I.branch[19].l_um_iw[159] ,
    \top_I.branch[19].l_um_iw[158] ,
    \top_I.branch[19].l_um_iw[157] ,
    \top_I.branch[19].l_um_iw[156] ,
    \top_I.branch[19].l_um_iw[155] ,
    \top_I.branch[19].l_um_iw[154] ,
    \top_I.branch[19].l_um_iw[153] ,
    \top_I.branch[19].l_um_iw[152] ,
    \top_I.branch[19].l_um_iw[151] ,
    \top_I.branch[19].l_um_iw[150] ,
    \top_I.branch[19].l_um_iw[149] ,
    \top_I.branch[19].l_um_iw[148] ,
    \top_I.branch[19].l_um_iw[147] ,
    \top_I.branch[19].l_um_iw[146] ,
    \top_I.branch[19].l_um_iw[145] ,
    \top_I.branch[19].l_um_iw[144] ,
    \top_I.branch[19].l_um_iw[143] ,
    \top_I.branch[19].l_um_iw[142] ,
    \top_I.branch[19].l_um_iw[141] ,
    \top_I.branch[19].l_um_iw[140] ,
    \top_I.branch[19].l_um_iw[139] ,
    \top_I.branch[19].l_um_iw[138] ,
    \top_I.branch[19].l_um_iw[137] ,
    \top_I.branch[19].l_um_iw[136] ,
    \top_I.branch[19].l_um_iw[135] ,
    \top_I.branch[19].l_um_iw[134] ,
    \top_I.branch[19].l_um_iw[133] ,
    \top_I.branch[19].l_um_iw[132] ,
    \top_I.branch[19].l_um_iw[131] ,
    \top_I.branch[19].l_um_iw[130] ,
    \top_I.branch[19].l_um_iw[129] ,
    \top_I.branch[19].l_um_iw[128] ,
    \top_I.branch[19].l_um_iw[127] ,
    \top_I.branch[19].l_um_iw[126] ,
    \top_I.branch[19].l_um_iw[125] ,
    \top_I.branch[19].l_um_iw[124] ,
    \top_I.branch[19].l_um_iw[123] ,
    \top_I.branch[19].l_um_iw[122] ,
    \top_I.branch[19].l_um_iw[121] ,
    \top_I.branch[19].l_um_iw[120] ,
    \top_I.branch[19].l_um_iw[119] ,
    \top_I.branch[19].l_um_iw[118] ,
    \top_I.branch[19].l_um_iw[117] ,
    \top_I.branch[19].l_um_iw[116] ,
    \top_I.branch[19].l_um_iw[115] ,
    \top_I.branch[19].l_um_iw[114] ,
    \top_I.branch[19].l_um_iw[113] ,
    \top_I.branch[19].l_um_iw[112] ,
    \top_I.branch[19].l_um_iw[111] ,
    \top_I.branch[19].l_um_iw[110] ,
    \top_I.branch[19].l_um_iw[109] ,
    \top_I.branch[19].l_um_iw[108] ,
    \top_I.branch[19].l_um_iw[107] ,
    \top_I.branch[19].l_um_iw[106] ,
    \top_I.branch[19].l_um_iw[105] ,
    \top_I.branch[19].l_um_iw[104] ,
    \top_I.branch[19].l_um_iw[103] ,
    \top_I.branch[19].l_um_iw[102] ,
    \top_I.branch[19].l_um_iw[101] ,
    \top_I.branch[19].l_um_iw[100] ,
    \top_I.branch[19].l_um_iw[99] ,
    \top_I.branch[19].l_um_iw[98] ,
    \top_I.branch[19].l_um_iw[97] ,
    \top_I.branch[19].l_um_iw[96] ,
    \top_I.branch[19].l_um_iw[95] ,
    \top_I.branch[19].l_um_iw[94] ,
    \top_I.branch[19].l_um_iw[93] ,
    \top_I.branch[19].l_um_iw[92] ,
    \top_I.branch[19].l_um_iw[91] ,
    \top_I.branch[19].l_um_iw[90] ,
    \top_I.branch[19].l_um_iw[89] ,
    \top_I.branch[19].l_um_iw[88] ,
    \top_I.branch[19].l_um_iw[87] ,
    \top_I.branch[19].l_um_iw[86] ,
    \top_I.branch[19].l_um_iw[85] ,
    \top_I.branch[19].l_um_iw[84] ,
    \top_I.branch[19].l_um_iw[83] ,
    \top_I.branch[19].l_um_iw[82] ,
    \top_I.branch[19].l_um_iw[81] ,
    \top_I.branch[19].l_um_iw[80] ,
    \top_I.branch[19].l_um_iw[79] ,
    \top_I.branch[19].l_um_iw[78] ,
    \top_I.branch[19].l_um_iw[77] ,
    \top_I.branch[19].l_um_iw[76] ,
    \top_I.branch[19].l_um_iw[75] ,
    \top_I.branch[19].l_um_iw[74] ,
    \top_I.branch[19].l_um_iw[73] ,
    \top_I.branch[19].l_um_iw[72] ,
    \top_I.branch[19].l_um_iw[71] ,
    \top_I.branch[19].l_um_iw[70] ,
    \top_I.branch[19].l_um_iw[69] ,
    \top_I.branch[19].l_um_iw[68] ,
    \top_I.branch[19].l_um_iw[67] ,
    \top_I.branch[19].l_um_iw[66] ,
    \top_I.branch[19].l_um_iw[65] ,
    \top_I.branch[19].l_um_iw[64] ,
    \top_I.branch[19].l_um_iw[63] ,
    \top_I.branch[19].l_um_iw[62] ,
    \top_I.branch[19].l_um_iw[61] ,
    \top_I.branch[19].l_um_iw[60] ,
    \top_I.branch[19].l_um_iw[59] ,
    \top_I.branch[19].l_um_iw[58] ,
    \top_I.branch[19].l_um_iw[57] ,
    \top_I.branch[19].l_um_iw[56] ,
    \top_I.branch[19].l_um_iw[55] ,
    \top_I.branch[19].l_um_iw[54] ,
    \top_I.branch[19].l_um_iw[53] ,
    \top_I.branch[19].l_um_iw[52] ,
    \top_I.branch[19].l_um_iw[51] ,
    \top_I.branch[19].l_um_iw[50] ,
    \top_I.branch[19].l_um_iw[49] ,
    \top_I.branch[19].l_um_iw[48] ,
    \top_I.branch[19].l_um_iw[47] ,
    \top_I.branch[19].l_um_iw[46] ,
    \top_I.branch[19].l_um_iw[45] ,
    \top_I.branch[19].l_um_iw[44] ,
    \top_I.branch[19].l_um_iw[43] ,
    \top_I.branch[19].l_um_iw[42] ,
    \top_I.branch[19].l_um_iw[41] ,
    \top_I.branch[19].l_um_iw[40] ,
    \top_I.branch[19].l_um_iw[39] ,
    \top_I.branch[19].l_um_iw[38] ,
    \top_I.branch[19].l_um_iw[37] ,
    \top_I.branch[19].l_um_iw[36] ,
    \top_I.branch[19].l_um_iw[35] ,
    \top_I.branch[19].l_um_iw[34] ,
    \top_I.branch[19].l_um_iw[33] ,
    \top_I.branch[19].l_um_iw[32] ,
    \top_I.branch[19].l_um_iw[31] ,
    \top_I.branch[19].l_um_iw[30] ,
    \top_I.branch[19].l_um_iw[29] ,
    \top_I.branch[19].l_um_iw[28] ,
    \top_I.branch[19].l_um_iw[27] ,
    \top_I.branch[19].l_um_iw[26] ,
    \top_I.branch[19].l_um_iw[25] ,
    \top_I.branch[19].l_um_iw[24] ,
    \top_I.branch[19].l_um_iw[23] ,
    \top_I.branch[19].l_um_iw[22] ,
    \top_I.branch[19].l_um_iw[21] ,
    \top_I.branch[19].l_um_iw[20] ,
    \top_I.branch[19].l_um_iw[19] ,
    \top_I.branch[19].l_um_iw[18] ,
    \top_I.branch[19].l_um_iw[17] ,
    \top_I.branch[19].l_um_iw[16] ,
    \top_I.branch[19].l_um_iw[15] ,
    \top_I.branch[19].l_um_iw[14] ,
    \top_I.branch[19].l_um_iw[13] ,
    \top_I.branch[19].l_um_iw[12] ,
    \top_I.branch[19].l_um_iw[11] ,
    \top_I.branch[19].l_um_iw[10] ,
    \top_I.branch[19].l_um_iw[9] ,
    \top_I.branch[19].l_um_iw[8] ,
    \top_I.branch[19].l_um_iw[7] ,
    \top_I.branch[19].l_um_iw[6] ,
    \top_I.branch[19].l_um_iw[5] ,
    \top_I.branch[19].l_um_iw[4] ,
    \top_I.branch[19].l_um_iw[3] ,
    \top_I.branch[19].l_um_iw[2] ,
    \top_I.branch[19].l_um_iw[1] ,
    \top_I.branch[19].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[1] ,
    \top_I.branch[19].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[15] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[14] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[13] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[12] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[11] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[10] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[9] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[8] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[7] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[6] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[5] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[4] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[3] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].l_um_k_zero[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[19].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] ,
    \top_I.branch[19].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[1].col_um[0].um_bot_I.block_0_16.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[0] ),
    .ena(\top_I.branch[1].l_um_ena[0] ),
    .rst_n(\top_I.branch[1].l_um_iw[1] ),
    .ui_in({\top_I.branch[1].l_um_iw[9] ,
    \top_I.branch[1].l_um_iw[8] ,
    \top_I.branch[1].l_um_iw[7] ,
    \top_I.branch[1].l_um_iw[6] ,
    \top_I.branch[1].l_um_iw[5] ,
    \top_I.branch[1].l_um_iw[4] ,
    \top_I.branch[1].l_um_iw[3] ,
    \top_I.branch[1].l_um_iw[2] }),
    .uio_in({\top_I.branch[1].l_um_iw[17] ,
    \top_I.branch[1].l_um_iw[16] ,
    \top_I.branch[1].l_um_iw[15] ,
    \top_I.branch[1].l_um_iw[14] ,
    \top_I.branch[1].l_um_iw[13] ,
    \top_I.branch[1].l_um_iw[12] ,
    \top_I.branch[1].l_um_iw[11] ,
    \top_I.branch[1].l_um_iw[10] }),
    .uio_oe({\top_I.branch[1].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_tomkeddie_a \top_I.branch[1].col_um[0].um_top_I.block_1_16.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[18] ),
    .ena(\top_I.branch[1].l_um_ena[1] ),
    .rst_n(\top_I.branch[1].l_um_iw[19] ),
    .ui_in({\top_I.branch[1].l_um_iw[27] ,
    \top_I.branch[1].l_um_iw[26] ,
    \top_I.branch[1].l_um_iw[25] ,
    \top_I.branch[1].l_um_iw[24] ,
    \top_I.branch[1].l_um_iw[23] ,
    \top_I.branch[1].l_um_iw[22] ,
    \top_I.branch[1].l_um_iw[21] ,
    \top_I.branch[1].l_um_iw[20] }),
    .uio_in({\top_I.branch[1].l_um_iw[35] ,
    \top_I.branch[1].l_um_iw[34] ,
    \top_I.branch[1].l_um_iw[33] ,
    \top_I.branch[1].l_um_iw[32] ,
    \top_I.branch[1].l_um_iw[31] ,
    \top_I.branch[1].l_um_iw[30] ,
    \top_I.branch[1].l_um_iw[29] ,
    \top_I.branch[1].l_um_iw[28] }),
    .uio_oe({\top_I.branch[1].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[0] }));
 tt_um_algofoogle_solo_squash \top_I.branch[1].col_um[1].um_bot_I.block_0_17.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[36] ),
    .ena(\top_I.branch[1].l_um_ena[2] ),
    .rst_n(\top_I.branch[1].l_um_iw[37] ),
    .ui_in({\top_I.branch[1].l_um_iw[45] ,
    \top_I.branch[1].l_um_iw[44] ,
    \top_I.branch[1].l_um_iw[43] ,
    \top_I.branch[1].l_um_iw[42] ,
    \top_I.branch[1].l_um_iw[41] ,
    \top_I.branch[1].l_um_iw[40] ,
    \top_I.branch[1].l_um_iw[39] ,
    \top_I.branch[1].l_um_iw[38] }),
    .uio_in({\top_I.branch[1].l_um_iw[53] ,
    \top_I.branch[1].l_um_iw[52] ,
    \top_I.branch[1].l_um_iw[51] ,
    \top_I.branch[1].l_um_iw[50] ,
    \top_I.branch[1].l_um_iw[49] ,
    \top_I.branch[1].l_um_iw[48] ,
    \top_I.branch[1].l_um_iw[47] ,
    \top_I.branch[1].l_um_iw[46] }),
    .uio_oe({\top_I.branch[1].col_um[1].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[1].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[1].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[0] }));
 tt_um_apu_pulse \top_I.branch[1].col_um[2].um_bot_I.block_0_18.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[72] ),
    .ena(\top_I.branch[1].l_um_ena[4] ),
    .rst_n(\top_I.branch[1].l_um_iw[73] ),
    .ui_in({\top_I.branch[1].l_um_iw[81] ,
    \top_I.branch[1].l_um_iw[80] ,
    \top_I.branch[1].l_um_iw[79] ,
    \top_I.branch[1].l_um_iw[78] ,
    \top_I.branch[1].l_um_iw[77] ,
    \top_I.branch[1].l_um_iw[76] ,
    \top_I.branch[1].l_um_iw[75] ,
    \top_I.branch[1].l_um_iw[74] }),
    .uio_in({\top_I.branch[1].l_um_iw[89] ,
    \top_I.branch[1].l_um_iw[88] ,
    \top_I.branch[1].l_um_iw[87] ,
    \top_I.branch[1].l_um_iw[86] ,
    \top_I.branch[1].l_um_iw[85] ,
    \top_I.branch[1].l_um_iw[84] ,
    \top_I.branch[1].l_um_iw[83] ,
    \top_I.branch[1].l_um_iw[82] }),
    .uio_oe({\top_I.branch[1].col_um[2].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[2].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[2].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[0] }));
 tt_um_htfab_totp \top_I.branch[1].col_um[2].um_top_I.block_1_18.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[90] ),
    .ena(\top_I.branch[1].l_um_ena[5] ),
    .rst_n(\top_I.branch[1].l_um_iw[91] ),
    .ui_in({\top_I.branch[1].l_um_iw[99] ,
    \top_I.branch[1].l_um_iw[98] ,
    \top_I.branch[1].l_um_iw[97] ,
    \top_I.branch[1].l_um_iw[96] ,
    \top_I.branch[1].l_um_iw[95] ,
    \top_I.branch[1].l_um_iw[94] ,
    \top_I.branch[1].l_um_iw[93] ,
    \top_I.branch[1].l_um_iw[92] }),
    .uio_in({\top_I.branch[1].l_um_iw[107] ,
    \top_I.branch[1].l_um_iw[106] ,
    \top_I.branch[1].l_um_iw[105] ,
    \top_I.branch[1].l_um_iw[104] ,
    \top_I.branch[1].l_um_iw[103] ,
    \top_I.branch[1].l_um_iw[102] ,
    \top_I.branch[1].l_um_iw[101] ,
    \top_I.branch[1].l_um_iw[100] }),
    .uio_oe({\top_I.branch[1].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[0] }));
 tt_um_thorkn_vgaclock \top_I.branch[1].col_um[3].um_bot_I.block_0_19.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[108] ),
    .ena(\top_I.branch[1].l_um_ena[6] ),
    .rst_n(\top_I.branch[1].l_um_iw[109] ),
    .ui_in({\top_I.branch[1].l_um_iw[117] ,
    \top_I.branch[1].l_um_iw[116] ,
    \top_I.branch[1].l_um_iw[115] ,
    \top_I.branch[1].l_um_iw[114] ,
    \top_I.branch[1].l_um_iw[113] ,
    \top_I.branch[1].l_um_iw[112] ,
    \top_I.branch[1].l_um_iw[111] ,
    \top_I.branch[1].l_um_iw[110] }),
    .uio_in({\top_I.branch[1].l_um_iw[125] ,
    \top_I.branch[1].l_um_iw[124] ,
    \top_I.branch[1].l_um_iw[123] ,
    \top_I.branch[1].l_um_iw[122] ,
    \top_I.branch[1].l_um_iw[121] ,
    \top_I.branch[1].l_um_iw[120] ,
    \top_I.branch[1].l_um_iw[119] ,
    \top_I.branch[1].l_um_iw[118] }),
    .uio_oe({\top_I.branch[1].col_um[3].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[3].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[3].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[0] }));
 tt_um_wokwi_347497504164545108 \top_I.branch[1].col_um[4].um_bot_I.block_0_20.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[144] ),
    .ena(\top_I.branch[1].l_um_ena[8] ),
    .rst_n(\top_I.branch[1].l_um_iw[145] ),
    .ui_in({\top_I.branch[1].l_um_iw[153] ,
    \top_I.branch[1].l_um_iw[152] ,
    \top_I.branch[1].l_um_iw[151] ,
    \top_I.branch[1].l_um_iw[150] ,
    \top_I.branch[1].l_um_iw[149] ,
    \top_I.branch[1].l_um_iw[148] ,
    \top_I.branch[1].l_um_iw[147] ,
    \top_I.branch[1].l_um_iw[146] }),
    .uio_in({\top_I.branch[1].l_um_iw[161] ,
    \top_I.branch[1].l_um_iw[160] ,
    \top_I.branch[1].l_um_iw[159] ,
    \top_I.branch[1].l_um_iw[158] ,
    \top_I.branch[1].l_um_iw[157] ,
    \top_I.branch[1].l_um_iw[156] ,
    \top_I.branch[1].l_um_iw[155] ,
    \top_I.branch[1].l_um_iw[154] }),
    .uio_oe({\top_I.branch[1].col_um[4].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[4].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[4].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[0] }));
 tt_um_Reloj_top \top_I.branch[1].col_um[4].um_top_I.block_1_20.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[162] ),
    .ena(\top_I.branch[1].l_um_ena[9] ),
    .rst_n(\top_I.branch[1].l_um_iw[163] ),
    .ui_in({\top_I.branch[1].l_um_iw[171] ,
    \top_I.branch[1].l_um_iw[170] ,
    \top_I.branch[1].l_um_iw[169] ,
    \top_I.branch[1].l_um_iw[168] ,
    \top_I.branch[1].l_um_iw[167] ,
    \top_I.branch[1].l_um_iw[166] ,
    \top_I.branch[1].l_um_iw[165] ,
    \top_I.branch[1].l_um_iw[164] }),
    .uio_in({\top_I.branch[1].l_um_iw[179] ,
    \top_I.branch[1].l_um_iw[178] ,
    \top_I.branch[1].l_um_iw[177] ,
    \top_I.branch[1].l_um_iw[176] ,
    \top_I.branch[1].l_um_iw[175] ,
    \top_I.branch[1].l_um_iw[174] ,
    \top_I.branch[1].l_um_iw[173] ,
    \top_I.branch[1].l_um_iw[172] }),
    .uio_oe({\top_I.branch[1].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[0] }));
 tt_um_wokwi_347144898258928211 \top_I.branch[1].col_um[5].um_bot_I.block_0_21.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[180] ),
    .ena(\top_I.branch[1].l_um_ena[10] ),
    .rst_n(\top_I.branch[1].l_um_iw[181] ),
    .ui_in({\top_I.branch[1].l_um_iw[189] ,
    \top_I.branch[1].l_um_iw[188] ,
    \top_I.branch[1].l_um_iw[187] ,
    \top_I.branch[1].l_um_iw[186] ,
    \top_I.branch[1].l_um_iw[185] ,
    \top_I.branch[1].l_um_iw[184] ,
    \top_I.branch[1].l_um_iw[183] ,
    \top_I.branch[1].l_um_iw[182] }),
    .uio_in({\top_I.branch[1].l_um_iw[197] ,
    \top_I.branch[1].l_um_iw[196] ,
    \top_I.branch[1].l_um_iw[195] ,
    \top_I.branch[1].l_um_iw[194] ,
    \top_I.branch[1].l_um_iw[193] ,
    \top_I.branch[1].l_um_iw[192] ,
    \top_I.branch[1].l_um_iw[191] ,
    \top_I.branch[1].l_um_iw[190] }),
    .uio_oe({\top_I.branch[1].col_um[5].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[5].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[5].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[0] }));
 tt_um_wokwi_347417602591556180 \top_I.branch[1].col_um[6].um_bot_I.block_0_22.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[216] ),
    .ena(\top_I.branch[1].l_um_ena[12] ),
    .rst_n(\top_I.branch[1].l_um_iw[217] ),
    .ui_in({\top_I.branch[1].l_um_iw[225] ,
    \top_I.branch[1].l_um_iw[224] ,
    \top_I.branch[1].l_um_iw[223] ,
    \top_I.branch[1].l_um_iw[222] ,
    \top_I.branch[1].l_um_iw[221] ,
    \top_I.branch[1].l_um_iw[220] ,
    \top_I.branch[1].l_um_iw[219] ,
    \top_I.branch[1].l_um_iw[218] }),
    .uio_in({\top_I.branch[1].l_um_iw[233] ,
    \top_I.branch[1].l_um_iw[232] ,
    \top_I.branch[1].l_um_iw[231] ,
    \top_I.branch[1].l_um_iw[230] ,
    \top_I.branch[1].l_um_iw[229] ,
    \top_I.branch[1].l_um_iw[228] ,
    \top_I.branch[1].l_um_iw[227] ,
    \top_I.branch[1].l_um_iw[226] }),
    .uio_oe({\top_I.branch[1].col_um[6].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[6].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[6].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[0] }));
 tt_um_urish_simon \top_I.branch[1].col_um[6].um_top_I.block_1_22.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[234] ),
    .ena(\top_I.branch[1].l_um_ena[13] ),
    .rst_n(\top_I.branch[1].l_um_iw[235] ),
    .ui_in({\top_I.branch[1].l_um_iw[243] ,
    \top_I.branch[1].l_um_iw[242] ,
    \top_I.branch[1].l_um_iw[241] ,
    \top_I.branch[1].l_um_iw[240] ,
    \top_I.branch[1].l_um_iw[239] ,
    \top_I.branch[1].l_um_iw[238] ,
    \top_I.branch[1].l_um_iw[237] ,
    \top_I.branch[1].l_um_iw[236] }),
    .uio_in({\top_I.branch[1].l_um_iw[251] ,
    \top_I.branch[1].l_um_iw[250] ,
    \top_I.branch[1].l_um_iw[249] ,
    \top_I.branch[1].l_um_iw[248] ,
    \top_I.branch[1].l_um_iw[247] ,
    \top_I.branch[1].l_um_iw[246] ,
    \top_I.branch[1].l_um_iw[245] ,
    \top_I.branch[1].l_um_iw[244] }),
    .uio_oe({\top_I.branch[1].col_um[6].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[6].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[6].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[0] }));
 tt_um_psychogenic_neptuneproportional \top_I.branch[1].col_um[7].um_bot_I.block_0_23.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[252] ),
    .ena(\top_I.branch[1].l_um_ena[14] ),
    .rst_n(\top_I.branch[1].l_um_iw[253] ),
    .ui_in({\top_I.branch[1].l_um_iw[261] ,
    \top_I.branch[1].l_um_iw[260] ,
    \top_I.branch[1].l_um_iw[259] ,
    \top_I.branch[1].l_um_iw[258] ,
    \top_I.branch[1].l_um_iw[257] ,
    \top_I.branch[1].l_um_iw[256] ,
    \top_I.branch[1].l_um_iw[255] ,
    \top_I.branch[1].l_um_iw[254] }),
    .uio_in({\top_I.branch[1].l_um_iw[269] ,
    \top_I.branch[1].l_um_iw[268] ,
    \top_I.branch[1].l_um_iw[267] ,
    \top_I.branch[1].l_um_iw[266] ,
    \top_I.branch[1].l_um_iw[265] ,
    \top_I.branch[1].l_um_iw[264] ,
    \top_I.branch[1].l_um_iw[263] ,
    \top_I.branch[1].l_um_iw[262] }),
    .uio_oe({\top_I.branch[1].col_um[7].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[7].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[7].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[0] }));
 tt_um_kiwih_tt_top \top_I.branch[1].col_um[7].um_top_I.block_1_23.tt_um_I  (.clk(\top_I.branch[1].l_um_iw[270] ),
    .ena(\top_I.branch[1].l_um_ena[15] ),
    .rst_n(\top_I.branch[1].l_um_iw[271] ),
    .ui_in({\top_I.branch[1].l_um_iw[279] ,
    \top_I.branch[1].l_um_iw[278] ,
    \top_I.branch[1].l_um_iw[277] ,
    \top_I.branch[1].l_um_iw[276] ,
    \top_I.branch[1].l_um_iw[275] ,
    \top_I.branch[1].l_um_iw[274] ,
    \top_I.branch[1].l_um_iw[273] ,
    \top_I.branch[1].l_um_iw[272] }),
    .uio_in({\top_I.branch[1].l_um_iw[287] ,
    \top_I.branch[1].l_um_iw[286] ,
    \top_I.branch[1].l_um_iw[285] ,
    \top_I.branch[1].l_um_iw[284] ,
    \top_I.branch[1].l_um_iw[283] ,
    \top_I.branch[1].l_um_iw[282] ,
    \top_I.branch[1].l_um_iw[281] ,
    \top_I.branch[1].l_um_iw[280] }),
    .uio_oe({\top_I.branch[1].col_um[7].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[1].col_um[7].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[1].col_um[7].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[1].mux_I  (.k_one(\top_I.branch[1].l_k_one ),
    .k_zero(\top_I.branch[1].l_k_zero ),
    .addr({\top_I.branch[1].l_k_zero ,
    \top_I.branch[1].l_k_zero ,
    \top_I.branch[1].l_k_zero ,
    \top_I.branch[1].l_k_zero ,
    \top_I.branch[1].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[1].l_um_ena[15] ,
    \top_I.branch[1].l_um_ena[14] ,
    \top_I.branch[1].l_um_ena[13] ,
    \top_I.branch[1].l_um_ena[12] ,
    \top_I.branch[1].l_um_ena[11] ,
    \top_I.branch[1].l_um_ena[10] ,
    \top_I.branch[1].l_um_ena[9] ,
    \top_I.branch[1].l_um_ena[8] ,
    \top_I.branch[1].l_um_ena[7] ,
    \top_I.branch[1].l_um_ena[6] ,
    \top_I.branch[1].l_um_ena[5] ,
    \top_I.branch[1].l_um_ena[4] ,
    \top_I.branch[1].l_um_ena[3] ,
    \top_I.branch[1].l_um_ena[2] ,
    \top_I.branch[1].l_um_ena[1] ,
    \top_I.branch[1].l_um_ena[0] }),
    .um_iw({\top_I.branch[1].l_um_iw[287] ,
    \top_I.branch[1].l_um_iw[286] ,
    \top_I.branch[1].l_um_iw[285] ,
    \top_I.branch[1].l_um_iw[284] ,
    \top_I.branch[1].l_um_iw[283] ,
    \top_I.branch[1].l_um_iw[282] ,
    \top_I.branch[1].l_um_iw[281] ,
    \top_I.branch[1].l_um_iw[280] ,
    \top_I.branch[1].l_um_iw[279] ,
    \top_I.branch[1].l_um_iw[278] ,
    \top_I.branch[1].l_um_iw[277] ,
    \top_I.branch[1].l_um_iw[276] ,
    \top_I.branch[1].l_um_iw[275] ,
    \top_I.branch[1].l_um_iw[274] ,
    \top_I.branch[1].l_um_iw[273] ,
    \top_I.branch[1].l_um_iw[272] ,
    \top_I.branch[1].l_um_iw[271] ,
    \top_I.branch[1].l_um_iw[270] ,
    \top_I.branch[1].l_um_iw[269] ,
    \top_I.branch[1].l_um_iw[268] ,
    \top_I.branch[1].l_um_iw[267] ,
    \top_I.branch[1].l_um_iw[266] ,
    \top_I.branch[1].l_um_iw[265] ,
    \top_I.branch[1].l_um_iw[264] ,
    \top_I.branch[1].l_um_iw[263] ,
    \top_I.branch[1].l_um_iw[262] ,
    \top_I.branch[1].l_um_iw[261] ,
    \top_I.branch[1].l_um_iw[260] ,
    \top_I.branch[1].l_um_iw[259] ,
    \top_I.branch[1].l_um_iw[258] ,
    \top_I.branch[1].l_um_iw[257] ,
    \top_I.branch[1].l_um_iw[256] ,
    \top_I.branch[1].l_um_iw[255] ,
    \top_I.branch[1].l_um_iw[254] ,
    \top_I.branch[1].l_um_iw[253] ,
    \top_I.branch[1].l_um_iw[252] ,
    \top_I.branch[1].l_um_iw[251] ,
    \top_I.branch[1].l_um_iw[250] ,
    \top_I.branch[1].l_um_iw[249] ,
    \top_I.branch[1].l_um_iw[248] ,
    \top_I.branch[1].l_um_iw[247] ,
    \top_I.branch[1].l_um_iw[246] ,
    \top_I.branch[1].l_um_iw[245] ,
    \top_I.branch[1].l_um_iw[244] ,
    \top_I.branch[1].l_um_iw[243] ,
    \top_I.branch[1].l_um_iw[242] ,
    \top_I.branch[1].l_um_iw[241] ,
    \top_I.branch[1].l_um_iw[240] ,
    \top_I.branch[1].l_um_iw[239] ,
    \top_I.branch[1].l_um_iw[238] ,
    \top_I.branch[1].l_um_iw[237] ,
    \top_I.branch[1].l_um_iw[236] ,
    \top_I.branch[1].l_um_iw[235] ,
    \top_I.branch[1].l_um_iw[234] ,
    \top_I.branch[1].l_um_iw[233] ,
    \top_I.branch[1].l_um_iw[232] ,
    \top_I.branch[1].l_um_iw[231] ,
    \top_I.branch[1].l_um_iw[230] ,
    \top_I.branch[1].l_um_iw[229] ,
    \top_I.branch[1].l_um_iw[228] ,
    \top_I.branch[1].l_um_iw[227] ,
    \top_I.branch[1].l_um_iw[226] ,
    \top_I.branch[1].l_um_iw[225] ,
    \top_I.branch[1].l_um_iw[224] ,
    \top_I.branch[1].l_um_iw[223] ,
    \top_I.branch[1].l_um_iw[222] ,
    \top_I.branch[1].l_um_iw[221] ,
    \top_I.branch[1].l_um_iw[220] ,
    \top_I.branch[1].l_um_iw[219] ,
    \top_I.branch[1].l_um_iw[218] ,
    \top_I.branch[1].l_um_iw[217] ,
    \top_I.branch[1].l_um_iw[216] ,
    \top_I.branch[1].l_um_iw[215] ,
    \top_I.branch[1].l_um_iw[214] ,
    \top_I.branch[1].l_um_iw[213] ,
    \top_I.branch[1].l_um_iw[212] ,
    \top_I.branch[1].l_um_iw[211] ,
    \top_I.branch[1].l_um_iw[210] ,
    \top_I.branch[1].l_um_iw[209] ,
    \top_I.branch[1].l_um_iw[208] ,
    \top_I.branch[1].l_um_iw[207] ,
    \top_I.branch[1].l_um_iw[206] ,
    \top_I.branch[1].l_um_iw[205] ,
    \top_I.branch[1].l_um_iw[204] ,
    \top_I.branch[1].l_um_iw[203] ,
    \top_I.branch[1].l_um_iw[202] ,
    \top_I.branch[1].l_um_iw[201] ,
    \top_I.branch[1].l_um_iw[200] ,
    \top_I.branch[1].l_um_iw[199] ,
    \top_I.branch[1].l_um_iw[198] ,
    \top_I.branch[1].l_um_iw[197] ,
    \top_I.branch[1].l_um_iw[196] ,
    \top_I.branch[1].l_um_iw[195] ,
    \top_I.branch[1].l_um_iw[194] ,
    \top_I.branch[1].l_um_iw[193] ,
    \top_I.branch[1].l_um_iw[192] ,
    \top_I.branch[1].l_um_iw[191] ,
    \top_I.branch[1].l_um_iw[190] ,
    \top_I.branch[1].l_um_iw[189] ,
    \top_I.branch[1].l_um_iw[188] ,
    \top_I.branch[1].l_um_iw[187] ,
    \top_I.branch[1].l_um_iw[186] ,
    \top_I.branch[1].l_um_iw[185] ,
    \top_I.branch[1].l_um_iw[184] ,
    \top_I.branch[1].l_um_iw[183] ,
    \top_I.branch[1].l_um_iw[182] ,
    \top_I.branch[1].l_um_iw[181] ,
    \top_I.branch[1].l_um_iw[180] ,
    \top_I.branch[1].l_um_iw[179] ,
    \top_I.branch[1].l_um_iw[178] ,
    \top_I.branch[1].l_um_iw[177] ,
    \top_I.branch[1].l_um_iw[176] ,
    \top_I.branch[1].l_um_iw[175] ,
    \top_I.branch[1].l_um_iw[174] ,
    \top_I.branch[1].l_um_iw[173] ,
    \top_I.branch[1].l_um_iw[172] ,
    \top_I.branch[1].l_um_iw[171] ,
    \top_I.branch[1].l_um_iw[170] ,
    \top_I.branch[1].l_um_iw[169] ,
    \top_I.branch[1].l_um_iw[168] ,
    \top_I.branch[1].l_um_iw[167] ,
    \top_I.branch[1].l_um_iw[166] ,
    \top_I.branch[1].l_um_iw[165] ,
    \top_I.branch[1].l_um_iw[164] ,
    \top_I.branch[1].l_um_iw[163] ,
    \top_I.branch[1].l_um_iw[162] ,
    \top_I.branch[1].l_um_iw[161] ,
    \top_I.branch[1].l_um_iw[160] ,
    \top_I.branch[1].l_um_iw[159] ,
    \top_I.branch[1].l_um_iw[158] ,
    \top_I.branch[1].l_um_iw[157] ,
    \top_I.branch[1].l_um_iw[156] ,
    \top_I.branch[1].l_um_iw[155] ,
    \top_I.branch[1].l_um_iw[154] ,
    \top_I.branch[1].l_um_iw[153] ,
    \top_I.branch[1].l_um_iw[152] ,
    \top_I.branch[1].l_um_iw[151] ,
    \top_I.branch[1].l_um_iw[150] ,
    \top_I.branch[1].l_um_iw[149] ,
    \top_I.branch[1].l_um_iw[148] ,
    \top_I.branch[1].l_um_iw[147] ,
    \top_I.branch[1].l_um_iw[146] ,
    \top_I.branch[1].l_um_iw[145] ,
    \top_I.branch[1].l_um_iw[144] ,
    \top_I.branch[1].l_um_iw[143] ,
    \top_I.branch[1].l_um_iw[142] ,
    \top_I.branch[1].l_um_iw[141] ,
    \top_I.branch[1].l_um_iw[140] ,
    \top_I.branch[1].l_um_iw[139] ,
    \top_I.branch[1].l_um_iw[138] ,
    \top_I.branch[1].l_um_iw[137] ,
    \top_I.branch[1].l_um_iw[136] ,
    \top_I.branch[1].l_um_iw[135] ,
    \top_I.branch[1].l_um_iw[134] ,
    \top_I.branch[1].l_um_iw[133] ,
    \top_I.branch[1].l_um_iw[132] ,
    \top_I.branch[1].l_um_iw[131] ,
    \top_I.branch[1].l_um_iw[130] ,
    \top_I.branch[1].l_um_iw[129] ,
    \top_I.branch[1].l_um_iw[128] ,
    \top_I.branch[1].l_um_iw[127] ,
    \top_I.branch[1].l_um_iw[126] ,
    \top_I.branch[1].l_um_iw[125] ,
    \top_I.branch[1].l_um_iw[124] ,
    \top_I.branch[1].l_um_iw[123] ,
    \top_I.branch[1].l_um_iw[122] ,
    \top_I.branch[1].l_um_iw[121] ,
    \top_I.branch[1].l_um_iw[120] ,
    \top_I.branch[1].l_um_iw[119] ,
    \top_I.branch[1].l_um_iw[118] ,
    \top_I.branch[1].l_um_iw[117] ,
    \top_I.branch[1].l_um_iw[116] ,
    \top_I.branch[1].l_um_iw[115] ,
    \top_I.branch[1].l_um_iw[114] ,
    \top_I.branch[1].l_um_iw[113] ,
    \top_I.branch[1].l_um_iw[112] ,
    \top_I.branch[1].l_um_iw[111] ,
    \top_I.branch[1].l_um_iw[110] ,
    \top_I.branch[1].l_um_iw[109] ,
    \top_I.branch[1].l_um_iw[108] ,
    \top_I.branch[1].l_um_iw[107] ,
    \top_I.branch[1].l_um_iw[106] ,
    \top_I.branch[1].l_um_iw[105] ,
    \top_I.branch[1].l_um_iw[104] ,
    \top_I.branch[1].l_um_iw[103] ,
    \top_I.branch[1].l_um_iw[102] ,
    \top_I.branch[1].l_um_iw[101] ,
    \top_I.branch[1].l_um_iw[100] ,
    \top_I.branch[1].l_um_iw[99] ,
    \top_I.branch[1].l_um_iw[98] ,
    \top_I.branch[1].l_um_iw[97] ,
    \top_I.branch[1].l_um_iw[96] ,
    \top_I.branch[1].l_um_iw[95] ,
    \top_I.branch[1].l_um_iw[94] ,
    \top_I.branch[1].l_um_iw[93] ,
    \top_I.branch[1].l_um_iw[92] ,
    \top_I.branch[1].l_um_iw[91] ,
    \top_I.branch[1].l_um_iw[90] ,
    \top_I.branch[1].l_um_iw[89] ,
    \top_I.branch[1].l_um_iw[88] ,
    \top_I.branch[1].l_um_iw[87] ,
    \top_I.branch[1].l_um_iw[86] ,
    \top_I.branch[1].l_um_iw[85] ,
    \top_I.branch[1].l_um_iw[84] ,
    \top_I.branch[1].l_um_iw[83] ,
    \top_I.branch[1].l_um_iw[82] ,
    \top_I.branch[1].l_um_iw[81] ,
    \top_I.branch[1].l_um_iw[80] ,
    \top_I.branch[1].l_um_iw[79] ,
    \top_I.branch[1].l_um_iw[78] ,
    \top_I.branch[1].l_um_iw[77] ,
    \top_I.branch[1].l_um_iw[76] ,
    \top_I.branch[1].l_um_iw[75] ,
    \top_I.branch[1].l_um_iw[74] ,
    \top_I.branch[1].l_um_iw[73] ,
    \top_I.branch[1].l_um_iw[72] ,
    \top_I.branch[1].l_um_iw[71] ,
    \top_I.branch[1].l_um_iw[70] ,
    \top_I.branch[1].l_um_iw[69] ,
    \top_I.branch[1].l_um_iw[68] ,
    \top_I.branch[1].l_um_iw[67] ,
    \top_I.branch[1].l_um_iw[66] ,
    \top_I.branch[1].l_um_iw[65] ,
    \top_I.branch[1].l_um_iw[64] ,
    \top_I.branch[1].l_um_iw[63] ,
    \top_I.branch[1].l_um_iw[62] ,
    \top_I.branch[1].l_um_iw[61] ,
    \top_I.branch[1].l_um_iw[60] ,
    \top_I.branch[1].l_um_iw[59] ,
    \top_I.branch[1].l_um_iw[58] ,
    \top_I.branch[1].l_um_iw[57] ,
    \top_I.branch[1].l_um_iw[56] ,
    \top_I.branch[1].l_um_iw[55] ,
    \top_I.branch[1].l_um_iw[54] ,
    \top_I.branch[1].l_um_iw[53] ,
    \top_I.branch[1].l_um_iw[52] ,
    \top_I.branch[1].l_um_iw[51] ,
    \top_I.branch[1].l_um_iw[50] ,
    \top_I.branch[1].l_um_iw[49] ,
    \top_I.branch[1].l_um_iw[48] ,
    \top_I.branch[1].l_um_iw[47] ,
    \top_I.branch[1].l_um_iw[46] ,
    \top_I.branch[1].l_um_iw[45] ,
    \top_I.branch[1].l_um_iw[44] ,
    \top_I.branch[1].l_um_iw[43] ,
    \top_I.branch[1].l_um_iw[42] ,
    \top_I.branch[1].l_um_iw[41] ,
    \top_I.branch[1].l_um_iw[40] ,
    \top_I.branch[1].l_um_iw[39] ,
    \top_I.branch[1].l_um_iw[38] ,
    \top_I.branch[1].l_um_iw[37] ,
    \top_I.branch[1].l_um_iw[36] ,
    \top_I.branch[1].l_um_iw[35] ,
    \top_I.branch[1].l_um_iw[34] ,
    \top_I.branch[1].l_um_iw[33] ,
    \top_I.branch[1].l_um_iw[32] ,
    \top_I.branch[1].l_um_iw[31] ,
    \top_I.branch[1].l_um_iw[30] ,
    \top_I.branch[1].l_um_iw[29] ,
    \top_I.branch[1].l_um_iw[28] ,
    \top_I.branch[1].l_um_iw[27] ,
    \top_I.branch[1].l_um_iw[26] ,
    \top_I.branch[1].l_um_iw[25] ,
    \top_I.branch[1].l_um_iw[24] ,
    \top_I.branch[1].l_um_iw[23] ,
    \top_I.branch[1].l_um_iw[22] ,
    \top_I.branch[1].l_um_iw[21] ,
    \top_I.branch[1].l_um_iw[20] ,
    \top_I.branch[1].l_um_iw[19] ,
    \top_I.branch[1].l_um_iw[18] ,
    \top_I.branch[1].l_um_iw[17] ,
    \top_I.branch[1].l_um_iw[16] ,
    \top_I.branch[1].l_um_iw[15] ,
    \top_I.branch[1].l_um_iw[14] ,
    \top_I.branch[1].l_um_iw[13] ,
    \top_I.branch[1].l_um_iw[12] ,
    \top_I.branch[1].l_um_iw[11] ,
    \top_I.branch[1].l_um_iw[10] ,
    \top_I.branch[1].l_um_iw[9] ,
    \top_I.branch[1].l_um_iw[8] ,
    \top_I.branch[1].l_um_iw[7] ,
    \top_I.branch[1].l_um_iw[6] ,
    \top_I.branch[1].l_um_iw[5] ,
    \top_I.branch[1].l_um_iw[4] ,
    \top_I.branch[1].l_um_iw[3] ,
    \top_I.branch[1].l_um_iw[2] ,
    \top_I.branch[1].l_um_iw[1] ,
    \top_I.branch[1].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[1].l_um_k_zero[15] ,
    \top_I.branch[1].l_um_k_zero[14] ,
    \top_I.branch[1].l_um_k_zero[13] ,
    \top_I.branch[1].l_um_k_zero[12] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[10] ,
    \top_I.branch[1].l_um_k_zero[9] ,
    \top_I.branch[1].l_um_k_zero[8] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[6] ,
    \top_I.branch[1].l_um_k_zero[5] ,
    \top_I.branch[1].l_um_k_zero[4] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[2] ,
    \top_I.branch[1].l_um_k_zero[1] ,
    \top_I.branch[1].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[1].col_um[7].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_oe[0] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uio_out[0] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[7].um_top_I.uo_out[0] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[7].um_bot_I.uo_out[0] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_oe[0] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uio_out[0] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[6].um_top_I.uo_out[0] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[6].um_bot_I.uo_out[0] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].l_um_k_zero[11] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[5].um_bot_I.uo_out[0] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_oe[0] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uio_out[0] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[4].um_top_I.uo_out[0] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[4].um_bot_I.uo_out[0] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].l_um_k_zero[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[3].um_bot_I.uo_out[0] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_oe[0] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uio_out[0] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[2].um_top_I.uo_out[0] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[2].um_bot_I.uo_out[0] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].l_um_k_zero[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[1].um_bot_I.uo_out[0] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[1].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[1].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[20].col_um[0].um_bot_I.block_20_0.tt_um_I  (.clk(\top_I.branch[20].l_um_iw[0] ),
    .ena(\top_I.branch[20].l_um_ena[0] ),
    .rst_n(\top_I.branch[20].l_um_iw[1] ),
    .ui_in({\top_I.branch[20].l_um_iw[9] ,
    \top_I.branch[20].l_um_iw[8] ,
    \top_I.branch[20].l_um_iw[7] ,
    \top_I.branch[20].l_um_iw[6] ,
    \top_I.branch[20].l_um_iw[5] ,
    \top_I.branch[20].l_um_iw[4] ,
    \top_I.branch[20].l_um_iw[3] ,
    \top_I.branch[20].l_um_iw[2] }),
    .uio_in({\top_I.branch[20].l_um_iw[17] ,
    \top_I.branch[20].l_um_iw[16] ,
    \top_I.branch[20].l_um_iw[15] ,
    \top_I.branch[20].l_um_iw[14] ,
    \top_I.branch[20].l_um_iw[13] ,
    \top_I.branch[20].l_um_iw[12] ,
    \top_I.branch[20].l_um_iw[11] ,
    \top_I.branch[20].l_um_iw[10] }),
    .uio_oe({\top_I.branch[20].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[20].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[20].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[20].mux_I  (.k_one(\top_I.branch[20].l_k_one ),
    .k_zero(\top_I.branch[20].l_k_zero ),
    .addr({\top_I.branch[20].l_k_one ,
    \top_I.branch[20].l_k_zero ,
    \top_I.branch[20].l_k_one ,
    \top_I.branch[20].l_k_zero ,
    \top_I.branch[20].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[20].l_um_ena[15] ,
    \top_I.branch[20].l_um_ena[14] ,
    \top_I.branch[20].l_um_ena[13] ,
    \top_I.branch[20].l_um_ena[12] ,
    \top_I.branch[20].l_um_ena[11] ,
    \top_I.branch[20].l_um_ena[10] ,
    \top_I.branch[20].l_um_ena[9] ,
    \top_I.branch[20].l_um_ena[8] ,
    \top_I.branch[20].l_um_ena[7] ,
    \top_I.branch[20].l_um_ena[6] ,
    \top_I.branch[20].l_um_ena[5] ,
    \top_I.branch[20].l_um_ena[4] ,
    \top_I.branch[20].l_um_ena[3] ,
    \top_I.branch[20].l_um_ena[2] ,
    \top_I.branch[20].l_um_ena[1] ,
    \top_I.branch[20].l_um_ena[0] }),
    .um_iw({\top_I.branch[20].l_um_iw[287] ,
    \top_I.branch[20].l_um_iw[286] ,
    \top_I.branch[20].l_um_iw[285] ,
    \top_I.branch[20].l_um_iw[284] ,
    \top_I.branch[20].l_um_iw[283] ,
    \top_I.branch[20].l_um_iw[282] ,
    \top_I.branch[20].l_um_iw[281] ,
    \top_I.branch[20].l_um_iw[280] ,
    \top_I.branch[20].l_um_iw[279] ,
    \top_I.branch[20].l_um_iw[278] ,
    \top_I.branch[20].l_um_iw[277] ,
    \top_I.branch[20].l_um_iw[276] ,
    \top_I.branch[20].l_um_iw[275] ,
    \top_I.branch[20].l_um_iw[274] ,
    \top_I.branch[20].l_um_iw[273] ,
    \top_I.branch[20].l_um_iw[272] ,
    \top_I.branch[20].l_um_iw[271] ,
    \top_I.branch[20].l_um_iw[270] ,
    \top_I.branch[20].l_um_iw[269] ,
    \top_I.branch[20].l_um_iw[268] ,
    \top_I.branch[20].l_um_iw[267] ,
    \top_I.branch[20].l_um_iw[266] ,
    \top_I.branch[20].l_um_iw[265] ,
    \top_I.branch[20].l_um_iw[264] ,
    \top_I.branch[20].l_um_iw[263] ,
    \top_I.branch[20].l_um_iw[262] ,
    \top_I.branch[20].l_um_iw[261] ,
    \top_I.branch[20].l_um_iw[260] ,
    \top_I.branch[20].l_um_iw[259] ,
    \top_I.branch[20].l_um_iw[258] ,
    \top_I.branch[20].l_um_iw[257] ,
    \top_I.branch[20].l_um_iw[256] ,
    \top_I.branch[20].l_um_iw[255] ,
    \top_I.branch[20].l_um_iw[254] ,
    \top_I.branch[20].l_um_iw[253] ,
    \top_I.branch[20].l_um_iw[252] ,
    \top_I.branch[20].l_um_iw[251] ,
    \top_I.branch[20].l_um_iw[250] ,
    \top_I.branch[20].l_um_iw[249] ,
    \top_I.branch[20].l_um_iw[248] ,
    \top_I.branch[20].l_um_iw[247] ,
    \top_I.branch[20].l_um_iw[246] ,
    \top_I.branch[20].l_um_iw[245] ,
    \top_I.branch[20].l_um_iw[244] ,
    \top_I.branch[20].l_um_iw[243] ,
    \top_I.branch[20].l_um_iw[242] ,
    \top_I.branch[20].l_um_iw[241] ,
    \top_I.branch[20].l_um_iw[240] ,
    \top_I.branch[20].l_um_iw[239] ,
    \top_I.branch[20].l_um_iw[238] ,
    \top_I.branch[20].l_um_iw[237] ,
    \top_I.branch[20].l_um_iw[236] ,
    \top_I.branch[20].l_um_iw[235] ,
    \top_I.branch[20].l_um_iw[234] ,
    \top_I.branch[20].l_um_iw[233] ,
    \top_I.branch[20].l_um_iw[232] ,
    \top_I.branch[20].l_um_iw[231] ,
    \top_I.branch[20].l_um_iw[230] ,
    \top_I.branch[20].l_um_iw[229] ,
    \top_I.branch[20].l_um_iw[228] ,
    \top_I.branch[20].l_um_iw[227] ,
    \top_I.branch[20].l_um_iw[226] ,
    \top_I.branch[20].l_um_iw[225] ,
    \top_I.branch[20].l_um_iw[224] ,
    \top_I.branch[20].l_um_iw[223] ,
    \top_I.branch[20].l_um_iw[222] ,
    \top_I.branch[20].l_um_iw[221] ,
    \top_I.branch[20].l_um_iw[220] ,
    \top_I.branch[20].l_um_iw[219] ,
    \top_I.branch[20].l_um_iw[218] ,
    \top_I.branch[20].l_um_iw[217] ,
    \top_I.branch[20].l_um_iw[216] ,
    \top_I.branch[20].l_um_iw[215] ,
    \top_I.branch[20].l_um_iw[214] ,
    \top_I.branch[20].l_um_iw[213] ,
    \top_I.branch[20].l_um_iw[212] ,
    \top_I.branch[20].l_um_iw[211] ,
    \top_I.branch[20].l_um_iw[210] ,
    \top_I.branch[20].l_um_iw[209] ,
    \top_I.branch[20].l_um_iw[208] ,
    \top_I.branch[20].l_um_iw[207] ,
    \top_I.branch[20].l_um_iw[206] ,
    \top_I.branch[20].l_um_iw[205] ,
    \top_I.branch[20].l_um_iw[204] ,
    \top_I.branch[20].l_um_iw[203] ,
    \top_I.branch[20].l_um_iw[202] ,
    \top_I.branch[20].l_um_iw[201] ,
    \top_I.branch[20].l_um_iw[200] ,
    \top_I.branch[20].l_um_iw[199] ,
    \top_I.branch[20].l_um_iw[198] ,
    \top_I.branch[20].l_um_iw[197] ,
    \top_I.branch[20].l_um_iw[196] ,
    \top_I.branch[20].l_um_iw[195] ,
    \top_I.branch[20].l_um_iw[194] ,
    \top_I.branch[20].l_um_iw[193] ,
    \top_I.branch[20].l_um_iw[192] ,
    \top_I.branch[20].l_um_iw[191] ,
    \top_I.branch[20].l_um_iw[190] ,
    \top_I.branch[20].l_um_iw[189] ,
    \top_I.branch[20].l_um_iw[188] ,
    \top_I.branch[20].l_um_iw[187] ,
    \top_I.branch[20].l_um_iw[186] ,
    \top_I.branch[20].l_um_iw[185] ,
    \top_I.branch[20].l_um_iw[184] ,
    \top_I.branch[20].l_um_iw[183] ,
    \top_I.branch[20].l_um_iw[182] ,
    \top_I.branch[20].l_um_iw[181] ,
    \top_I.branch[20].l_um_iw[180] ,
    \top_I.branch[20].l_um_iw[179] ,
    \top_I.branch[20].l_um_iw[178] ,
    \top_I.branch[20].l_um_iw[177] ,
    \top_I.branch[20].l_um_iw[176] ,
    \top_I.branch[20].l_um_iw[175] ,
    \top_I.branch[20].l_um_iw[174] ,
    \top_I.branch[20].l_um_iw[173] ,
    \top_I.branch[20].l_um_iw[172] ,
    \top_I.branch[20].l_um_iw[171] ,
    \top_I.branch[20].l_um_iw[170] ,
    \top_I.branch[20].l_um_iw[169] ,
    \top_I.branch[20].l_um_iw[168] ,
    \top_I.branch[20].l_um_iw[167] ,
    \top_I.branch[20].l_um_iw[166] ,
    \top_I.branch[20].l_um_iw[165] ,
    \top_I.branch[20].l_um_iw[164] ,
    \top_I.branch[20].l_um_iw[163] ,
    \top_I.branch[20].l_um_iw[162] ,
    \top_I.branch[20].l_um_iw[161] ,
    \top_I.branch[20].l_um_iw[160] ,
    \top_I.branch[20].l_um_iw[159] ,
    \top_I.branch[20].l_um_iw[158] ,
    \top_I.branch[20].l_um_iw[157] ,
    \top_I.branch[20].l_um_iw[156] ,
    \top_I.branch[20].l_um_iw[155] ,
    \top_I.branch[20].l_um_iw[154] ,
    \top_I.branch[20].l_um_iw[153] ,
    \top_I.branch[20].l_um_iw[152] ,
    \top_I.branch[20].l_um_iw[151] ,
    \top_I.branch[20].l_um_iw[150] ,
    \top_I.branch[20].l_um_iw[149] ,
    \top_I.branch[20].l_um_iw[148] ,
    \top_I.branch[20].l_um_iw[147] ,
    \top_I.branch[20].l_um_iw[146] ,
    \top_I.branch[20].l_um_iw[145] ,
    \top_I.branch[20].l_um_iw[144] ,
    \top_I.branch[20].l_um_iw[143] ,
    \top_I.branch[20].l_um_iw[142] ,
    \top_I.branch[20].l_um_iw[141] ,
    \top_I.branch[20].l_um_iw[140] ,
    \top_I.branch[20].l_um_iw[139] ,
    \top_I.branch[20].l_um_iw[138] ,
    \top_I.branch[20].l_um_iw[137] ,
    \top_I.branch[20].l_um_iw[136] ,
    \top_I.branch[20].l_um_iw[135] ,
    \top_I.branch[20].l_um_iw[134] ,
    \top_I.branch[20].l_um_iw[133] ,
    \top_I.branch[20].l_um_iw[132] ,
    \top_I.branch[20].l_um_iw[131] ,
    \top_I.branch[20].l_um_iw[130] ,
    \top_I.branch[20].l_um_iw[129] ,
    \top_I.branch[20].l_um_iw[128] ,
    \top_I.branch[20].l_um_iw[127] ,
    \top_I.branch[20].l_um_iw[126] ,
    \top_I.branch[20].l_um_iw[125] ,
    \top_I.branch[20].l_um_iw[124] ,
    \top_I.branch[20].l_um_iw[123] ,
    \top_I.branch[20].l_um_iw[122] ,
    \top_I.branch[20].l_um_iw[121] ,
    \top_I.branch[20].l_um_iw[120] ,
    \top_I.branch[20].l_um_iw[119] ,
    \top_I.branch[20].l_um_iw[118] ,
    \top_I.branch[20].l_um_iw[117] ,
    \top_I.branch[20].l_um_iw[116] ,
    \top_I.branch[20].l_um_iw[115] ,
    \top_I.branch[20].l_um_iw[114] ,
    \top_I.branch[20].l_um_iw[113] ,
    \top_I.branch[20].l_um_iw[112] ,
    \top_I.branch[20].l_um_iw[111] ,
    \top_I.branch[20].l_um_iw[110] ,
    \top_I.branch[20].l_um_iw[109] ,
    \top_I.branch[20].l_um_iw[108] ,
    \top_I.branch[20].l_um_iw[107] ,
    \top_I.branch[20].l_um_iw[106] ,
    \top_I.branch[20].l_um_iw[105] ,
    \top_I.branch[20].l_um_iw[104] ,
    \top_I.branch[20].l_um_iw[103] ,
    \top_I.branch[20].l_um_iw[102] ,
    \top_I.branch[20].l_um_iw[101] ,
    \top_I.branch[20].l_um_iw[100] ,
    \top_I.branch[20].l_um_iw[99] ,
    \top_I.branch[20].l_um_iw[98] ,
    \top_I.branch[20].l_um_iw[97] ,
    \top_I.branch[20].l_um_iw[96] ,
    \top_I.branch[20].l_um_iw[95] ,
    \top_I.branch[20].l_um_iw[94] ,
    \top_I.branch[20].l_um_iw[93] ,
    \top_I.branch[20].l_um_iw[92] ,
    \top_I.branch[20].l_um_iw[91] ,
    \top_I.branch[20].l_um_iw[90] ,
    \top_I.branch[20].l_um_iw[89] ,
    \top_I.branch[20].l_um_iw[88] ,
    \top_I.branch[20].l_um_iw[87] ,
    \top_I.branch[20].l_um_iw[86] ,
    \top_I.branch[20].l_um_iw[85] ,
    \top_I.branch[20].l_um_iw[84] ,
    \top_I.branch[20].l_um_iw[83] ,
    \top_I.branch[20].l_um_iw[82] ,
    \top_I.branch[20].l_um_iw[81] ,
    \top_I.branch[20].l_um_iw[80] ,
    \top_I.branch[20].l_um_iw[79] ,
    \top_I.branch[20].l_um_iw[78] ,
    \top_I.branch[20].l_um_iw[77] ,
    \top_I.branch[20].l_um_iw[76] ,
    \top_I.branch[20].l_um_iw[75] ,
    \top_I.branch[20].l_um_iw[74] ,
    \top_I.branch[20].l_um_iw[73] ,
    \top_I.branch[20].l_um_iw[72] ,
    \top_I.branch[20].l_um_iw[71] ,
    \top_I.branch[20].l_um_iw[70] ,
    \top_I.branch[20].l_um_iw[69] ,
    \top_I.branch[20].l_um_iw[68] ,
    \top_I.branch[20].l_um_iw[67] ,
    \top_I.branch[20].l_um_iw[66] ,
    \top_I.branch[20].l_um_iw[65] ,
    \top_I.branch[20].l_um_iw[64] ,
    \top_I.branch[20].l_um_iw[63] ,
    \top_I.branch[20].l_um_iw[62] ,
    \top_I.branch[20].l_um_iw[61] ,
    \top_I.branch[20].l_um_iw[60] ,
    \top_I.branch[20].l_um_iw[59] ,
    \top_I.branch[20].l_um_iw[58] ,
    \top_I.branch[20].l_um_iw[57] ,
    \top_I.branch[20].l_um_iw[56] ,
    \top_I.branch[20].l_um_iw[55] ,
    \top_I.branch[20].l_um_iw[54] ,
    \top_I.branch[20].l_um_iw[53] ,
    \top_I.branch[20].l_um_iw[52] ,
    \top_I.branch[20].l_um_iw[51] ,
    \top_I.branch[20].l_um_iw[50] ,
    \top_I.branch[20].l_um_iw[49] ,
    \top_I.branch[20].l_um_iw[48] ,
    \top_I.branch[20].l_um_iw[47] ,
    \top_I.branch[20].l_um_iw[46] ,
    \top_I.branch[20].l_um_iw[45] ,
    \top_I.branch[20].l_um_iw[44] ,
    \top_I.branch[20].l_um_iw[43] ,
    \top_I.branch[20].l_um_iw[42] ,
    \top_I.branch[20].l_um_iw[41] ,
    \top_I.branch[20].l_um_iw[40] ,
    \top_I.branch[20].l_um_iw[39] ,
    \top_I.branch[20].l_um_iw[38] ,
    \top_I.branch[20].l_um_iw[37] ,
    \top_I.branch[20].l_um_iw[36] ,
    \top_I.branch[20].l_um_iw[35] ,
    \top_I.branch[20].l_um_iw[34] ,
    \top_I.branch[20].l_um_iw[33] ,
    \top_I.branch[20].l_um_iw[32] ,
    \top_I.branch[20].l_um_iw[31] ,
    \top_I.branch[20].l_um_iw[30] ,
    \top_I.branch[20].l_um_iw[29] ,
    \top_I.branch[20].l_um_iw[28] ,
    \top_I.branch[20].l_um_iw[27] ,
    \top_I.branch[20].l_um_iw[26] ,
    \top_I.branch[20].l_um_iw[25] ,
    \top_I.branch[20].l_um_iw[24] ,
    \top_I.branch[20].l_um_iw[23] ,
    \top_I.branch[20].l_um_iw[22] ,
    \top_I.branch[20].l_um_iw[21] ,
    \top_I.branch[20].l_um_iw[20] ,
    \top_I.branch[20].l_um_iw[19] ,
    \top_I.branch[20].l_um_iw[18] ,
    \top_I.branch[20].l_um_iw[17] ,
    \top_I.branch[20].l_um_iw[16] ,
    \top_I.branch[20].l_um_iw[15] ,
    \top_I.branch[20].l_um_iw[14] ,
    \top_I.branch[20].l_um_iw[13] ,
    \top_I.branch[20].l_um_iw[12] ,
    \top_I.branch[20].l_um_iw[11] ,
    \top_I.branch[20].l_um_iw[10] ,
    \top_I.branch[20].l_um_iw[9] ,
    \top_I.branch[20].l_um_iw[8] ,
    \top_I.branch[20].l_um_iw[7] ,
    \top_I.branch[20].l_um_iw[6] ,
    \top_I.branch[20].l_um_iw[5] ,
    \top_I.branch[20].l_um_iw[4] ,
    \top_I.branch[20].l_um_iw[3] ,
    \top_I.branch[20].l_um_iw[2] ,
    \top_I.branch[20].l_um_iw[1] ,
    \top_I.branch[20].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[15] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[14] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[13] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[12] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[11] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[10] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[9] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[8] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[7] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[6] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[5] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[4] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[3] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[2] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].l_um_k_zero[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[20].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[21].col_um[0].um_bot_I.block_20_16.tt_um_I  (.clk(\top_I.branch[21].l_um_iw[0] ),
    .ena(\top_I.branch[21].l_um_ena[0] ),
    .rst_n(\top_I.branch[21].l_um_iw[1] ),
    .ui_in({\top_I.branch[21].l_um_iw[9] ,
    \top_I.branch[21].l_um_iw[8] ,
    \top_I.branch[21].l_um_iw[7] ,
    \top_I.branch[21].l_um_iw[6] ,
    \top_I.branch[21].l_um_iw[5] ,
    \top_I.branch[21].l_um_iw[4] ,
    \top_I.branch[21].l_um_iw[3] ,
    \top_I.branch[21].l_um_iw[2] }),
    .uio_in({\top_I.branch[21].l_um_iw[17] ,
    \top_I.branch[21].l_um_iw[16] ,
    \top_I.branch[21].l_um_iw[15] ,
    \top_I.branch[21].l_um_iw[14] ,
    \top_I.branch[21].l_um_iw[13] ,
    \top_I.branch[21].l_um_iw[12] ,
    \top_I.branch[21].l_um_iw[11] ,
    \top_I.branch[21].l_um_iw[10] }),
    .uio_oe({\top_I.branch[21].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[21].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[21].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[21].mux_I  (.k_one(\top_I.branch[21].l_k_one ),
    .k_zero(\top_I.branch[21].l_k_zero ),
    .addr({\top_I.branch[21].l_k_one ,
    \top_I.branch[21].l_k_zero ,
    \top_I.branch[21].l_k_one ,
    \top_I.branch[21].l_k_zero ,
    \top_I.branch[21].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[21].l_um_ena[15] ,
    \top_I.branch[21].l_um_ena[14] ,
    \top_I.branch[21].l_um_ena[13] ,
    \top_I.branch[21].l_um_ena[12] ,
    \top_I.branch[21].l_um_ena[11] ,
    \top_I.branch[21].l_um_ena[10] ,
    \top_I.branch[21].l_um_ena[9] ,
    \top_I.branch[21].l_um_ena[8] ,
    \top_I.branch[21].l_um_ena[7] ,
    \top_I.branch[21].l_um_ena[6] ,
    \top_I.branch[21].l_um_ena[5] ,
    \top_I.branch[21].l_um_ena[4] ,
    \top_I.branch[21].l_um_ena[3] ,
    \top_I.branch[21].l_um_ena[2] ,
    \top_I.branch[21].l_um_ena[1] ,
    \top_I.branch[21].l_um_ena[0] }),
    .um_iw({\top_I.branch[21].l_um_iw[287] ,
    \top_I.branch[21].l_um_iw[286] ,
    \top_I.branch[21].l_um_iw[285] ,
    \top_I.branch[21].l_um_iw[284] ,
    \top_I.branch[21].l_um_iw[283] ,
    \top_I.branch[21].l_um_iw[282] ,
    \top_I.branch[21].l_um_iw[281] ,
    \top_I.branch[21].l_um_iw[280] ,
    \top_I.branch[21].l_um_iw[279] ,
    \top_I.branch[21].l_um_iw[278] ,
    \top_I.branch[21].l_um_iw[277] ,
    \top_I.branch[21].l_um_iw[276] ,
    \top_I.branch[21].l_um_iw[275] ,
    \top_I.branch[21].l_um_iw[274] ,
    \top_I.branch[21].l_um_iw[273] ,
    \top_I.branch[21].l_um_iw[272] ,
    \top_I.branch[21].l_um_iw[271] ,
    \top_I.branch[21].l_um_iw[270] ,
    \top_I.branch[21].l_um_iw[269] ,
    \top_I.branch[21].l_um_iw[268] ,
    \top_I.branch[21].l_um_iw[267] ,
    \top_I.branch[21].l_um_iw[266] ,
    \top_I.branch[21].l_um_iw[265] ,
    \top_I.branch[21].l_um_iw[264] ,
    \top_I.branch[21].l_um_iw[263] ,
    \top_I.branch[21].l_um_iw[262] ,
    \top_I.branch[21].l_um_iw[261] ,
    \top_I.branch[21].l_um_iw[260] ,
    \top_I.branch[21].l_um_iw[259] ,
    \top_I.branch[21].l_um_iw[258] ,
    \top_I.branch[21].l_um_iw[257] ,
    \top_I.branch[21].l_um_iw[256] ,
    \top_I.branch[21].l_um_iw[255] ,
    \top_I.branch[21].l_um_iw[254] ,
    \top_I.branch[21].l_um_iw[253] ,
    \top_I.branch[21].l_um_iw[252] ,
    \top_I.branch[21].l_um_iw[251] ,
    \top_I.branch[21].l_um_iw[250] ,
    \top_I.branch[21].l_um_iw[249] ,
    \top_I.branch[21].l_um_iw[248] ,
    \top_I.branch[21].l_um_iw[247] ,
    \top_I.branch[21].l_um_iw[246] ,
    \top_I.branch[21].l_um_iw[245] ,
    \top_I.branch[21].l_um_iw[244] ,
    \top_I.branch[21].l_um_iw[243] ,
    \top_I.branch[21].l_um_iw[242] ,
    \top_I.branch[21].l_um_iw[241] ,
    \top_I.branch[21].l_um_iw[240] ,
    \top_I.branch[21].l_um_iw[239] ,
    \top_I.branch[21].l_um_iw[238] ,
    \top_I.branch[21].l_um_iw[237] ,
    \top_I.branch[21].l_um_iw[236] ,
    \top_I.branch[21].l_um_iw[235] ,
    \top_I.branch[21].l_um_iw[234] ,
    \top_I.branch[21].l_um_iw[233] ,
    \top_I.branch[21].l_um_iw[232] ,
    \top_I.branch[21].l_um_iw[231] ,
    \top_I.branch[21].l_um_iw[230] ,
    \top_I.branch[21].l_um_iw[229] ,
    \top_I.branch[21].l_um_iw[228] ,
    \top_I.branch[21].l_um_iw[227] ,
    \top_I.branch[21].l_um_iw[226] ,
    \top_I.branch[21].l_um_iw[225] ,
    \top_I.branch[21].l_um_iw[224] ,
    \top_I.branch[21].l_um_iw[223] ,
    \top_I.branch[21].l_um_iw[222] ,
    \top_I.branch[21].l_um_iw[221] ,
    \top_I.branch[21].l_um_iw[220] ,
    \top_I.branch[21].l_um_iw[219] ,
    \top_I.branch[21].l_um_iw[218] ,
    \top_I.branch[21].l_um_iw[217] ,
    \top_I.branch[21].l_um_iw[216] ,
    \top_I.branch[21].l_um_iw[215] ,
    \top_I.branch[21].l_um_iw[214] ,
    \top_I.branch[21].l_um_iw[213] ,
    \top_I.branch[21].l_um_iw[212] ,
    \top_I.branch[21].l_um_iw[211] ,
    \top_I.branch[21].l_um_iw[210] ,
    \top_I.branch[21].l_um_iw[209] ,
    \top_I.branch[21].l_um_iw[208] ,
    \top_I.branch[21].l_um_iw[207] ,
    \top_I.branch[21].l_um_iw[206] ,
    \top_I.branch[21].l_um_iw[205] ,
    \top_I.branch[21].l_um_iw[204] ,
    \top_I.branch[21].l_um_iw[203] ,
    \top_I.branch[21].l_um_iw[202] ,
    \top_I.branch[21].l_um_iw[201] ,
    \top_I.branch[21].l_um_iw[200] ,
    \top_I.branch[21].l_um_iw[199] ,
    \top_I.branch[21].l_um_iw[198] ,
    \top_I.branch[21].l_um_iw[197] ,
    \top_I.branch[21].l_um_iw[196] ,
    \top_I.branch[21].l_um_iw[195] ,
    \top_I.branch[21].l_um_iw[194] ,
    \top_I.branch[21].l_um_iw[193] ,
    \top_I.branch[21].l_um_iw[192] ,
    \top_I.branch[21].l_um_iw[191] ,
    \top_I.branch[21].l_um_iw[190] ,
    \top_I.branch[21].l_um_iw[189] ,
    \top_I.branch[21].l_um_iw[188] ,
    \top_I.branch[21].l_um_iw[187] ,
    \top_I.branch[21].l_um_iw[186] ,
    \top_I.branch[21].l_um_iw[185] ,
    \top_I.branch[21].l_um_iw[184] ,
    \top_I.branch[21].l_um_iw[183] ,
    \top_I.branch[21].l_um_iw[182] ,
    \top_I.branch[21].l_um_iw[181] ,
    \top_I.branch[21].l_um_iw[180] ,
    \top_I.branch[21].l_um_iw[179] ,
    \top_I.branch[21].l_um_iw[178] ,
    \top_I.branch[21].l_um_iw[177] ,
    \top_I.branch[21].l_um_iw[176] ,
    \top_I.branch[21].l_um_iw[175] ,
    \top_I.branch[21].l_um_iw[174] ,
    \top_I.branch[21].l_um_iw[173] ,
    \top_I.branch[21].l_um_iw[172] ,
    \top_I.branch[21].l_um_iw[171] ,
    \top_I.branch[21].l_um_iw[170] ,
    \top_I.branch[21].l_um_iw[169] ,
    \top_I.branch[21].l_um_iw[168] ,
    \top_I.branch[21].l_um_iw[167] ,
    \top_I.branch[21].l_um_iw[166] ,
    \top_I.branch[21].l_um_iw[165] ,
    \top_I.branch[21].l_um_iw[164] ,
    \top_I.branch[21].l_um_iw[163] ,
    \top_I.branch[21].l_um_iw[162] ,
    \top_I.branch[21].l_um_iw[161] ,
    \top_I.branch[21].l_um_iw[160] ,
    \top_I.branch[21].l_um_iw[159] ,
    \top_I.branch[21].l_um_iw[158] ,
    \top_I.branch[21].l_um_iw[157] ,
    \top_I.branch[21].l_um_iw[156] ,
    \top_I.branch[21].l_um_iw[155] ,
    \top_I.branch[21].l_um_iw[154] ,
    \top_I.branch[21].l_um_iw[153] ,
    \top_I.branch[21].l_um_iw[152] ,
    \top_I.branch[21].l_um_iw[151] ,
    \top_I.branch[21].l_um_iw[150] ,
    \top_I.branch[21].l_um_iw[149] ,
    \top_I.branch[21].l_um_iw[148] ,
    \top_I.branch[21].l_um_iw[147] ,
    \top_I.branch[21].l_um_iw[146] ,
    \top_I.branch[21].l_um_iw[145] ,
    \top_I.branch[21].l_um_iw[144] ,
    \top_I.branch[21].l_um_iw[143] ,
    \top_I.branch[21].l_um_iw[142] ,
    \top_I.branch[21].l_um_iw[141] ,
    \top_I.branch[21].l_um_iw[140] ,
    \top_I.branch[21].l_um_iw[139] ,
    \top_I.branch[21].l_um_iw[138] ,
    \top_I.branch[21].l_um_iw[137] ,
    \top_I.branch[21].l_um_iw[136] ,
    \top_I.branch[21].l_um_iw[135] ,
    \top_I.branch[21].l_um_iw[134] ,
    \top_I.branch[21].l_um_iw[133] ,
    \top_I.branch[21].l_um_iw[132] ,
    \top_I.branch[21].l_um_iw[131] ,
    \top_I.branch[21].l_um_iw[130] ,
    \top_I.branch[21].l_um_iw[129] ,
    \top_I.branch[21].l_um_iw[128] ,
    \top_I.branch[21].l_um_iw[127] ,
    \top_I.branch[21].l_um_iw[126] ,
    \top_I.branch[21].l_um_iw[125] ,
    \top_I.branch[21].l_um_iw[124] ,
    \top_I.branch[21].l_um_iw[123] ,
    \top_I.branch[21].l_um_iw[122] ,
    \top_I.branch[21].l_um_iw[121] ,
    \top_I.branch[21].l_um_iw[120] ,
    \top_I.branch[21].l_um_iw[119] ,
    \top_I.branch[21].l_um_iw[118] ,
    \top_I.branch[21].l_um_iw[117] ,
    \top_I.branch[21].l_um_iw[116] ,
    \top_I.branch[21].l_um_iw[115] ,
    \top_I.branch[21].l_um_iw[114] ,
    \top_I.branch[21].l_um_iw[113] ,
    \top_I.branch[21].l_um_iw[112] ,
    \top_I.branch[21].l_um_iw[111] ,
    \top_I.branch[21].l_um_iw[110] ,
    \top_I.branch[21].l_um_iw[109] ,
    \top_I.branch[21].l_um_iw[108] ,
    \top_I.branch[21].l_um_iw[107] ,
    \top_I.branch[21].l_um_iw[106] ,
    \top_I.branch[21].l_um_iw[105] ,
    \top_I.branch[21].l_um_iw[104] ,
    \top_I.branch[21].l_um_iw[103] ,
    \top_I.branch[21].l_um_iw[102] ,
    \top_I.branch[21].l_um_iw[101] ,
    \top_I.branch[21].l_um_iw[100] ,
    \top_I.branch[21].l_um_iw[99] ,
    \top_I.branch[21].l_um_iw[98] ,
    \top_I.branch[21].l_um_iw[97] ,
    \top_I.branch[21].l_um_iw[96] ,
    \top_I.branch[21].l_um_iw[95] ,
    \top_I.branch[21].l_um_iw[94] ,
    \top_I.branch[21].l_um_iw[93] ,
    \top_I.branch[21].l_um_iw[92] ,
    \top_I.branch[21].l_um_iw[91] ,
    \top_I.branch[21].l_um_iw[90] ,
    \top_I.branch[21].l_um_iw[89] ,
    \top_I.branch[21].l_um_iw[88] ,
    \top_I.branch[21].l_um_iw[87] ,
    \top_I.branch[21].l_um_iw[86] ,
    \top_I.branch[21].l_um_iw[85] ,
    \top_I.branch[21].l_um_iw[84] ,
    \top_I.branch[21].l_um_iw[83] ,
    \top_I.branch[21].l_um_iw[82] ,
    \top_I.branch[21].l_um_iw[81] ,
    \top_I.branch[21].l_um_iw[80] ,
    \top_I.branch[21].l_um_iw[79] ,
    \top_I.branch[21].l_um_iw[78] ,
    \top_I.branch[21].l_um_iw[77] ,
    \top_I.branch[21].l_um_iw[76] ,
    \top_I.branch[21].l_um_iw[75] ,
    \top_I.branch[21].l_um_iw[74] ,
    \top_I.branch[21].l_um_iw[73] ,
    \top_I.branch[21].l_um_iw[72] ,
    \top_I.branch[21].l_um_iw[71] ,
    \top_I.branch[21].l_um_iw[70] ,
    \top_I.branch[21].l_um_iw[69] ,
    \top_I.branch[21].l_um_iw[68] ,
    \top_I.branch[21].l_um_iw[67] ,
    \top_I.branch[21].l_um_iw[66] ,
    \top_I.branch[21].l_um_iw[65] ,
    \top_I.branch[21].l_um_iw[64] ,
    \top_I.branch[21].l_um_iw[63] ,
    \top_I.branch[21].l_um_iw[62] ,
    \top_I.branch[21].l_um_iw[61] ,
    \top_I.branch[21].l_um_iw[60] ,
    \top_I.branch[21].l_um_iw[59] ,
    \top_I.branch[21].l_um_iw[58] ,
    \top_I.branch[21].l_um_iw[57] ,
    \top_I.branch[21].l_um_iw[56] ,
    \top_I.branch[21].l_um_iw[55] ,
    \top_I.branch[21].l_um_iw[54] ,
    \top_I.branch[21].l_um_iw[53] ,
    \top_I.branch[21].l_um_iw[52] ,
    \top_I.branch[21].l_um_iw[51] ,
    \top_I.branch[21].l_um_iw[50] ,
    \top_I.branch[21].l_um_iw[49] ,
    \top_I.branch[21].l_um_iw[48] ,
    \top_I.branch[21].l_um_iw[47] ,
    \top_I.branch[21].l_um_iw[46] ,
    \top_I.branch[21].l_um_iw[45] ,
    \top_I.branch[21].l_um_iw[44] ,
    \top_I.branch[21].l_um_iw[43] ,
    \top_I.branch[21].l_um_iw[42] ,
    \top_I.branch[21].l_um_iw[41] ,
    \top_I.branch[21].l_um_iw[40] ,
    \top_I.branch[21].l_um_iw[39] ,
    \top_I.branch[21].l_um_iw[38] ,
    \top_I.branch[21].l_um_iw[37] ,
    \top_I.branch[21].l_um_iw[36] ,
    \top_I.branch[21].l_um_iw[35] ,
    \top_I.branch[21].l_um_iw[34] ,
    \top_I.branch[21].l_um_iw[33] ,
    \top_I.branch[21].l_um_iw[32] ,
    \top_I.branch[21].l_um_iw[31] ,
    \top_I.branch[21].l_um_iw[30] ,
    \top_I.branch[21].l_um_iw[29] ,
    \top_I.branch[21].l_um_iw[28] ,
    \top_I.branch[21].l_um_iw[27] ,
    \top_I.branch[21].l_um_iw[26] ,
    \top_I.branch[21].l_um_iw[25] ,
    \top_I.branch[21].l_um_iw[24] ,
    \top_I.branch[21].l_um_iw[23] ,
    \top_I.branch[21].l_um_iw[22] ,
    \top_I.branch[21].l_um_iw[21] ,
    \top_I.branch[21].l_um_iw[20] ,
    \top_I.branch[21].l_um_iw[19] ,
    \top_I.branch[21].l_um_iw[18] ,
    \top_I.branch[21].l_um_iw[17] ,
    \top_I.branch[21].l_um_iw[16] ,
    \top_I.branch[21].l_um_iw[15] ,
    \top_I.branch[21].l_um_iw[14] ,
    \top_I.branch[21].l_um_iw[13] ,
    \top_I.branch[21].l_um_iw[12] ,
    \top_I.branch[21].l_um_iw[11] ,
    \top_I.branch[21].l_um_iw[10] ,
    \top_I.branch[21].l_um_iw[9] ,
    \top_I.branch[21].l_um_iw[8] ,
    \top_I.branch[21].l_um_iw[7] ,
    \top_I.branch[21].l_um_iw[6] ,
    \top_I.branch[21].l_um_iw[5] ,
    \top_I.branch[21].l_um_iw[4] ,
    \top_I.branch[21].l_um_iw[3] ,
    \top_I.branch[21].l_um_iw[2] ,
    \top_I.branch[21].l_um_iw[1] ,
    \top_I.branch[21].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[15] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[14] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[13] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[12] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[11] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[10] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[9] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[8] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[7] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[6] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[5] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[4] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[3] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[2] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].l_um_k_zero[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[21].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[22].col_um[0].um_top_I.block_23_0.tt_um_I  (.clk(\top_I.branch[22].l_um_iw[18] ),
    .ena(\top_I.branch[22].l_um_ena[1] ),
    .rst_n(\top_I.branch[22].l_um_iw[19] ),
    .ui_in({\top_I.branch[22].l_um_iw[27] ,
    \top_I.branch[22].l_um_iw[26] ,
    \top_I.branch[22].l_um_iw[25] ,
    \top_I.branch[22].l_um_iw[24] ,
    \top_I.branch[22].l_um_iw[23] ,
    \top_I.branch[22].l_um_iw[22] ,
    \top_I.branch[22].l_um_iw[21] ,
    \top_I.branch[22].l_um_iw[20] }),
    .uio_in({\top_I.branch[22].l_um_iw[35] ,
    \top_I.branch[22].l_um_iw[34] ,
    \top_I.branch[22].l_um_iw[33] ,
    \top_I.branch[22].l_um_iw[32] ,
    \top_I.branch[22].l_um_iw[31] ,
    \top_I.branch[22].l_um_iw[30] ,
    \top_I.branch[22].l_um_iw[29] ,
    \top_I.branch[22].l_um_iw[28] }),
    .uio_oe({\top_I.branch[22].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[22].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[22].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[22].mux_I  (.k_one(\top_I.branch[22].l_k_one ),
    .k_zero(\top_I.branch[22].l_k_zero ),
    .addr({\top_I.branch[22].l_k_one ,
    \top_I.branch[22].l_k_zero ,
    \top_I.branch[22].l_k_one ,
    \top_I.branch[22].l_k_one ,
    \top_I.branch[22].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[22].l_um_ena[15] ,
    \top_I.branch[22].l_um_ena[14] ,
    \top_I.branch[22].l_um_ena[13] ,
    \top_I.branch[22].l_um_ena[12] ,
    \top_I.branch[22].l_um_ena[11] ,
    \top_I.branch[22].l_um_ena[10] ,
    \top_I.branch[22].l_um_ena[9] ,
    \top_I.branch[22].l_um_ena[8] ,
    \top_I.branch[22].l_um_ena[7] ,
    \top_I.branch[22].l_um_ena[6] ,
    \top_I.branch[22].l_um_ena[5] ,
    \top_I.branch[22].l_um_ena[4] ,
    \top_I.branch[22].l_um_ena[3] ,
    \top_I.branch[22].l_um_ena[2] ,
    \top_I.branch[22].l_um_ena[1] ,
    \top_I.branch[22].l_um_ena[0] }),
    .um_iw({\top_I.branch[22].l_um_iw[287] ,
    \top_I.branch[22].l_um_iw[286] ,
    \top_I.branch[22].l_um_iw[285] ,
    \top_I.branch[22].l_um_iw[284] ,
    \top_I.branch[22].l_um_iw[283] ,
    \top_I.branch[22].l_um_iw[282] ,
    \top_I.branch[22].l_um_iw[281] ,
    \top_I.branch[22].l_um_iw[280] ,
    \top_I.branch[22].l_um_iw[279] ,
    \top_I.branch[22].l_um_iw[278] ,
    \top_I.branch[22].l_um_iw[277] ,
    \top_I.branch[22].l_um_iw[276] ,
    \top_I.branch[22].l_um_iw[275] ,
    \top_I.branch[22].l_um_iw[274] ,
    \top_I.branch[22].l_um_iw[273] ,
    \top_I.branch[22].l_um_iw[272] ,
    \top_I.branch[22].l_um_iw[271] ,
    \top_I.branch[22].l_um_iw[270] ,
    \top_I.branch[22].l_um_iw[269] ,
    \top_I.branch[22].l_um_iw[268] ,
    \top_I.branch[22].l_um_iw[267] ,
    \top_I.branch[22].l_um_iw[266] ,
    \top_I.branch[22].l_um_iw[265] ,
    \top_I.branch[22].l_um_iw[264] ,
    \top_I.branch[22].l_um_iw[263] ,
    \top_I.branch[22].l_um_iw[262] ,
    \top_I.branch[22].l_um_iw[261] ,
    \top_I.branch[22].l_um_iw[260] ,
    \top_I.branch[22].l_um_iw[259] ,
    \top_I.branch[22].l_um_iw[258] ,
    \top_I.branch[22].l_um_iw[257] ,
    \top_I.branch[22].l_um_iw[256] ,
    \top_I.branch[22].l_um_iw[255] ,
    \top_I.branch[22].l_um_iw[254] ,
    \top_I.branch[22].l_um_iw[253] ,
    \top_I.branch[22].l_um_iw[252] ,
    \top_I.branch[22].l_um_iw[251] ,
    \top_I.branch[22].l_um_iw[250] ,
    \top_I.branch[22].l_um_iw[249] ,
    \top_I.branch[22].l_um_iw[248] ,
    \top_I.branch[22].l_um_iw[247] ,
    \top_I.branch[22].l_um_iw[246] ,
    \top_I.branch[22].l_um_iw[245] ,
    \top_I.branch[22].l_um_iw[244] ,
    \top_I.branch[22].l_um_iw[243] ,
    \top_I.branch[22].l_um_iw[242] ,
    \top_I.branch[22].l_um_iw[241] ,
    \top_I.branch[22].l_um_iw[240] ,
    \top_I.branch[22].l_um_iw[239] ,
    \top_I.branch[22].l_um_iw[238] ,
    \top_I.branch[22].l_um_iw[237] ,
    \top_I.branch[22].l_um_iw[236] ,
    \top_I.branch[22].l_um_iw[235] ,
    \top_I.branch[22].l_um_iw[234] ,
    \top_I.branch[22].l_um_iw[233] ,
    \top_I.branch[22].l_um_iw[232] ,
    \top_I.branch[22].l_um_iw[231] ,
    \top_I.branch[22].l_um_iw[230] ,
    \top_I.branch[22].l_um_iw[229] ,
    \top_I.branch[22].l_um_iw[228] ,
    \top_I.branch[22].l_um_iw[227] ,
    \top_I.branch[22].l_um_iw[226] ,
    \top_I.branch[22].l_um_iw[225] ,
    \top_I.branch[22].l_um_iw[224] ,
    \top_I.branch[22].l_um_iw[223] ,
    \top_I.branch[22].l_um_iw[222] ,
    \top_I.branch[22].l_um_iw[221] ,
    \top_I.branch[22].l_um_iw[220] ,
    \top_I.branch[22].l_um_iw[219] ,
    \top_I.branch[22].l_um_iw[218] ,
    \top_I.branch[22].l_um_iw[217] ,
    \top_I.branch[22].l_um_iw[216] ,
    \top_I.branch[22].l_um_iw[215] ,
    \top_I.branch[22].l_um_iw[214] ,
    \top_I.branch[22].l_um_iw[213] ,
    \top_I.branch[22].l_um_iw[212] ,
    \top_I.branch[22].l_um_iw[211] ,
    \top_I.branch[22].l_um_iw[210] ,
    \top_I.branch[22].l_um_iw[209] ,
    \top_I.branch[22].l_um_iw[208] ,
    \top_I.branch[22].l_um_iw[207] ,
    \top_I.branch[22].l_um_iw[206] ,
    \top_I.branch[22].l_um_iw[205] ,
    \top_I.branch[22].l_um_iw[204] ,
    \top_I.branch[22].l_um_iw[203] ,
    \top_I.branch[22].l_um_iw[202] ,
    \top_I.branch[22].l_um_iw[201] ,
    \top_I.branch[22].l_um_iw[200] ,
    \top_I.branch[22].l_um_iw[199] ,
    \top_I.branch[22].l_um_iw[198] ,
    \top_I.branch[22].l_um_iw[197] ,
    \top_I.branch[22].l_um_iw[196] ,
    \top_I.branch[22].l_um_iw[195] ,
    \top_I.branch[22].l_um_iw[194] ,
    \top_I.branch[22].l_um_iw[193] ,
    \top_I.branch[22].l_um_iw[192] ,
    \top_I.branch[22].l_um_iw[191] ,
    \top_I.branch[22].l_um_iw[190] ,
    \top_I.branch[22].l_um_iw[189] ,
    \top_I.branch[22].l_um_iw[188] ,
    \top_I.branch[22].l_um_iw[187] ,
    \top_I.branch[22].l_um_iw[186] ,
    \top_I.branch[22].l_um_iw[185] ,
    \top_I.branch[22].l_um_iw[184] ,
    \top_I.branch[22].l_um_iw[183] ,
    \top_I.branch[22].l_um_iw[182] ,
    \top_I.branch[22].l_um_iw[181] ,
    \top_I.branch[22].l_um_iw[180] ,
    \top_I.branch[22].l_um_iw[179] ,
    \top_I.branch[22].l_um_iw[178] ,
    \top_I.branch[22].l_um_iw[177] ,
    \top_I.branch[22].l_um_iw[176] ,
    \top_I.branch[22].l_um_iw[175] ,
    \top_I.branch[22].l_um_iw[174] ,
    \top_I.branch[22].l_um_iw[173] ,
    \top_I.branch[22].l_um_iw[172] ,
    \top_I.branch[22].l_um_iw[171] ,
    \top_I.branch[22].l_um_iw[170] ,
    \top_I.branch[22].l_um_iw[169] ,
    \top_I.branch[22].l_um_iw[168] ,
    \top_I.branch[22].l_um_iw[167] ,
    \top_I.branch[22].l_um_iw[166] ,
    \top_I.branch[22].l_um_iw[165] ,
    \top_I.branch[22].l_um_iw[164] ,
    \top_I.branch[22].l_um_iw[163] ,
    \top_I.branch[22].l_um_iw[162] ,
    \top_I.branch[22].l_um_iw[161] ,
    \top_I.branch[22].l_um_iw[160] ,
    \top_I.branch[22].l_um_iw[159] ,
    \top_I.branch[22].l_um_iw[158] ,
    \top_I.branch[22].l_um_iw[157] ,
    \top_I.branch[22].l_um_iw[156] ,
    \top_I.branch[22].l_um_iw[155] ,
    \top_I.branch[22].l_um_iw[154] ,
    \top_I.branch[22].l_um_iw[153] ,
    \top_I.branch[22].l_um_iw[152] ,
    \top_I.branch[22].l_um_iw[151] ,
    \top_I.branch[22].l_um_iw[150] ,
    \top_I.branch[22].l_um_iw[149] ,
    \top_I.branch[22].l_um_iw[148] ,
    \top_I.branch[22].l_um_iw[147] ,
    \top_I.branch[22].l_um_iw[146] ,
    \top_I.branch[22].l_um_iw[145] ,
    \top_I.branch[22].l_um_iw[144] ,
    \top_I.branch[22].l_um_iw[143] ,
    \top_I.branch[22].l_um_iw[142] ,
    \top_I.branch[22].l_um_iw[141] ,
    \top_I.branch[22].l_um_iw[140] ,
    \top_I.branch[22].l_um_iw[139] ,
    \top_I.branch[22].l_um_iw[138] ,
    \top_I.branch[22].l_um_iw[137] ,
    \top_I.branch[22].l_um_iw[136] ,
    \top_I.branch[22].l_um_iw[135] ,
    \top_I.branch[22].l_um_iw[134] ,
    \top_I.branch[22].l_um_iw[133] ,
    \top_I.branch[22].l_um_iw[132] ,
    \top_I.branch[22].l_um_iw[131] ,
    \top_I.branch[22].l_um_iw[130] ,
    \top_I.branch[22].l_um_iw[129] ,
    \top_I.branch[22].l_um_iw[128] ,
    \top_I.branch[22].l_um_iw[127] ,
    \top_I.branch[22].l_um_iw[126] ,
    \top_I.branch[22].l_um_iw[125] ,
    \top_I.branch[22].l_um_iw[124] ,
    \top_I.branch[22].l_um_iw[123] ,
    \top_I.branch[22].l_um_iw[122] ,
    \top_I.branch[22].l_um_iw[121] ,
    \top_I.branch[22].l_um_iw[120] ,
    \top_I.branch[22].l_um_iw[119] ,
    \top_I.branch[22].l_um_iw[118] ,
    \top_I.branch[22].l_um_iw[117] ,
    \top_I.branch[22].l_um_iw[116] ,
    \top_I.branch[22].l_um_iw[115] ,
    \top_I.branch[22].l_um_iw[114] ,
    \top_I.branch[22].l_um_iw[113] ,
    \top_I.branch[22].l_um_iw[112] ,
    \top_I.branch[22].l_um_iw[111] ,
    \top_I.branch[22].l_um_iw[110] ,
    \top_I.branch[22].l_um_iw[109] ,
    \top_I.branch[22].l_um_iw[108] ,
    \top_I.branch[22].l_um_iw[107] ,
    \top_I.branch[22].l_um_iw[106] ,
    \top_I.branch[22].l_um_iw[105] ,
    \top_I.branch[22].l_um_iw[104] ,
    \top_I.branch[22].l_um_iw[103] ,
    \top_I.branch[22].l_um_iw[102] ,
    \top_I.branch[22].l_um_iw[101] ,
    \top_I.branch[22].l_um_iw[100] ,
    \top_I.branch[22].l_um_iw[99] ,
    \top_I.branch[22].l_um_iw[98] ,
    \top_I.branch[22].l_um_iw[97] ,
    \top_I.branch[22].l_um_iw[96] ,
    \top_I.branch[22].l_um_iw[95] ,
    \top_I.branch[22].l_um_iw[94] ,
    \top_I.branch[22].l_um_iw[93] ,
    \top_I.branch[22].l_um_iw[92] ,
    \top_I.branch[22].l_um_iw[91] ,
    \top_I.branch[22].l_um_iw[90] ,
    \top_I.branch[22].l_um_iw[89] ,
    \top_I.branch[22].l_um_iw[88] ,
    \top_I.branch[22].l_um_iw[87] ,
    \top_I.branch[22].l_um_iw[86] ,
    \top_I.branch[22].l_um_iw[85] ,
    \top_I.branch[22].l_um_iw[84] ,
    \top_I.branch[22].l_um_iw[83] ,
    \top_I.branch[22].l_um_iw[82] ,
    \top_I.branch[22].l_um_iw[81] ,
    \top_I.branch[22].l_um_iw[80] ,
    \top_I.branch[22].l_um_iw[79] ,
    \top_I.branch[22].l_um_iw[78] ,
    \top_I.branch[22].l_um_iw[77] ,
    \top_I.branch[22].l_um_iw[76] ,
    \top_I.branch[22].l_um_iw[75] ,
    \top_I.branch[22].l_um_iw[74] ,
    \top_I.branch[22].l_um_iw[73] ,
    \top_I.branch[22].l_um_iw[72] ,
    \top_I.branch[22].l_um_iw[71] ,
    \top_I.branch[22].l_um_iw[70] ,
    \top_I.branch[22].l_um_iw[69] ,
    \top_I.branch[22].l_um_iw[68] ,
    \top_I.branch[22].l_um_iw[67] ,
    \top_I.branch[22].l_um_iw[66] ,
    \top_I.branch[22].l_um_iw[65] ,
    \top_I.branch[22].l_um_iw[64] ,
    \top_I.branch[22].l_um_iw[63] ,
    \top_I.branch[22].l_um_iw[62] ,
    \top_I.branch[22].l_um_iw[61] ,
    \top_I.branch[22].l_um_iw[60] ,
    \top_I.branch[22].l_um_iw[59] ,
    \top_I.branch[22].l_um_iw[58] ,
    \top_I.branch[22].l_um_iw[57] ,
    \top_I.branch[22].l_um_iw[56] ,
    \top_I.branch[22].l_um_iw[55] ,
    \top_I.branch[22].l_um_iw[54] ,
    \top_I.branch[22].l_um_iw[53] ,
    \top_I.branch[22].l_um_iw[52] ,
    \top_I.branch[22].l_um_iw[51] ,
    \top_I.branch[22].l_um_iw[50] ,
    \top_I.branch[22].l_um_iw[49] ,
    \top_I.branch[22].l_um_iw[48] ,
    \top_I.branch[22].l_um_iw[47] ,
    \top_I.branch[22].l_um_iw[46] ,
    \top_I.branch[22].l_um_iw[45] ,
    \top_I.branch[22].l_um_iw[44] ,
    \top_I.branch[22].l_um_iw[43] ,
    \top_I.branch[22].l_um_iw[42] ,
    \top_I.branch[22].l_um_iw[41] ,
    \top_I.branch[22].l_um_iw[40] ,
    \top_I.branch[22].l_um_iw[39] ,
    \top_I.branch[22].l_um_iw[38] ,
    \top_I.branch[22].l_um_iw[37] ,
    \top_I.branch[22].l_um_iw[36] ,
    \top_I.branch[22].l_um_iw[35] ,
    \top_I.branch[22].l_um_iw[34] ,
    \top_I.branch[22].l_um_iw[33] ,
    \top_I.branch[22].l_um_iw[32] ,
    \top_I.branch[22].l_um_iw[31] ,
    \top_I.branch[22].l_um_iw[30] ,
    \top_I.branch[22].l_um_iw[29] ,
    \top_I.branch[22].l_um_iw[28] ,
    \top_I.branch[22].l_um_iw[27] ,
    \top_I.branch[22].l_um_iw[26] ,
    \top_I.branch[22].l_um_iw[25] ,
    \top_I.branch[22].l_um_iw[24] ,
    \top_I.branch[22].l_um_iw[23] ,
    \top_I.branch[22].l_um_iw[22] ,
    \top_I.branch[22].l_um_iw[21] ,
    \top_I.branch[22].l_um_iw[20] ,
    \top_I.branch[22].l_um_iw[19] ,
    \top_I.branch[22].l_um_iw[18] ,
    \top_I.branch[22].l_um_iw[17] ,
    \top_I.branch[22].l_um_iw[16] ,
    \top_I.branch[22].l_um_iw[15] ,
    \top_I.branch[22].l_um_iw[14] ,
    \top_I.branch[22].l_um_iw[13] ,
    \top_I.branch[22].l_um_iw[12] ,
    \top_I.branch[22].l_um_iw[11] ,
    \top_I.branch[22].l_um_iw[10] ,
    \top_I.branch[22].l_um_iw[9] ,
    \top_I.branch[22].l_um_iw[8] ,
    \top_I.branch[22].l_um_iw[7] ,
    \top_I.branch[22].l_um_iw[6] ,
    \top_I.branch[22].l_um_iw[5] ,
    \top_I.branch[22].l_um_iw[4] ,
    \top_I.branch[22].l_um_iw[3] ,
    \top_I.branch[22].l_um_iw[2] ,
    \top_I.branch[22].l_um_iw[1] ,
    \top_I.branch[22].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[1] ,
    \top_I.branch[22].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[15] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[14] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[13] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[12] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[11] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[10] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[9] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[8] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[7] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[6] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[5] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[4] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[3] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].l_um_k_zero[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[22].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] ,
    \top_I.branch[22].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[23].col_um[0].um_top_I.block_23_16.tt_um_I  (.clk(\top_I.branch[23].l_um_iw[18] ),
    .ena(\top_I.branch[23].l_um_ena[1] ),
    .rst_n(\top_I.branch[23].l_um_iw[19] ),
    .ui_in({\top_I.branch[23].l_um_iw[27] ,
    \top_I.branch[23].l_um_iw[26] ,
    \top_I.branch[23].l_um_iw[25] ,
    \top_I.branch[23].l_um_iw[24] ,
    \top_I.branch[23].l_um_iw[23] ,
    \top_I.branch[23].l_um_iw[22] ,
    \top_I.branch[23].l_um_iw[21] ,
    \top_I.branch[23].l_um_iw[20] }),
    .uio_in({\top_I.branch[23].l_um_iw[35] ,
    \top_I.branch[23].l_um_iw[34] ,
    \top_I.branch[23].l_um_iw[33] ,
    \top_I.branch[23].l_um_iw[32] ,
    \top_I.branch[23].l_um_iw[31] ,
    \top_I.branch[23].l_um_iw[30] ,
    \top_I.branch[23].l_um_iw[29] ,
    \top_I.branch[23].l_um_iw[28] }),
    .uio_oe({\top_I.branch[23].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[23].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[23].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[23].mux_I  (.k_one(\top_I.branch[23].l_k_one ),
    .k_zero(\top_I.branch[23].l_k_zero ),
    .addr({\top_I.branch[23].l_k_one ,
    \top_I.branch[23].l_k_zero ,
    \top_I.branch[23].l_k_one ,
    \top_I.branch[23].l_k_one ,
    \top_I.branch[23].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[23].l_um_ena[15] ,
    \top_I.branch[23].l_um_ena[14] ,
    \top_I.branch[23].l_um_ena[13] ,
    \top_I.branch[23].l_um_ena[12] ,
    \top_I.branch[23].l_um_ena[11] ,
    \top_I.branch[23].l_um_ena[10] ,
    \top_I.branch[23].l_um_ena[9] ,
    \top_I.branch[23].l_um_ena[8] ,
    \top_I.branch[23].l_um_ena[7] ,
    \top_I.branch[23].l_um_ena[6] ,
    \top_I.branch[23].l_um_ena[5] ,
    \top_I.branch[23].l_um_ena[4] ,
    \top_I.branch[23].l_um_ena[3] ,
    \top_I.branch[23].l_um_ena[2] ,
    \top_I.branch[23].l_um_ena[1] ,
    \top_I.branch[23].l_um_ena[0] }),
    .um_iw({\top_I.branch[23].l_um_iw[287] ,
    \top_I.branch[23].l_um_iw[286] ,
    \top_I.branch[23].l_um_iw[285] ,
    \top_I.branch[23].l_um_iw[284] ,
    \top_I.branch[23].l_um_iw[283] ,
    \top_I.branch[23].l_um_iw[282] ,
    \top_I.branch[23].l_um_iw[281] ,
    \top_I.branch[23].l_um_iw[280] ,
    \top_I.branch[23].l_um_iw[279] ,
    \top_I.branch[23].l_um_iw[278] ,
    \top_I.branch[23].l_um_iw[277] ,
    \top_I.branch[23].l_um_iw[276] ,
    \top_I.branch[23].l_um_iw[275] ,
    \top_I.branch[23].l_um_iw[274] ,
    \top_I.branch[23].l_um_iw[273] ,
    \top_I.branch[23].l_um_iw[272] ,
    \top_I.branch[23].l_um_iw[271] ,
    \top_I.branch[23].l_um_iw[270] ,
    \top_I.branch[23].l_um_iw[269] ,
    \top_I.branch[23].l_um_iw[268] ,
    \top_I.branch[23].l_um_iw[267] ,
    \top_I.branch[23].l_um_iw[266] ,
    \top_I.branch[23].l_um_iw[265] ,
    \top_I.branch[23].l_um_iw[264] ,
    \top_I.branch[23].l_um_iw[263] ,
    \top_I.branch[23].l_um_iw[262] ,
    \top_I.branch[23].l_um_iw[261] ,
    \top_I.branch[23].l_um_iw[260] ,
    \top_I.branch[23].l_um_iw[259] ,
    \top_I.branch[23].l_um_iw[258] ,
    \top_I.branch[23].l_um_iw[257] ,
    \top_I.branch[23].l_um_iw[256] ,
    \top_I.branch[23].l_um_iw[255] ,
    \top_I.branch[23].l_um_iw[254] ,
    \top_I.branch[23].l_um_iw[253] ,
    \top_I.branch[23].l_um_iw[252] ,
    \top_I.branch[23].l_um_iw[251] ,
    \top_I.branch[23].l_um_iw[250] ,
    \top_I.branch[23].l_um_iw[249] ,
    \top_I.branch[23].l_um_iw[248] ,
    \top_I.branch[23].l_um_iw[247] ,
    \top_I.branch[23].l_um_iw[246] ,
    \top_I.branch[23].l_um_iw[245] ,
    \top_I.branch[23].l_um_iw[244] ,
    \top_I.branch[23].l_um_iw[243] ,
    \top_I.branch[23].l_um_iw[242] ,
    \top_I.branch[23].l_um_iw[241] ,
    \top_I.branch[23].l_um_iw[240] ,
    \top_I.branch[23].l_um_iw[239] ,
    \top_I.branch[23].l_um_iw[238] ,
    \top_I.branch[23].l_um_iw[237] ,
    \top_I.branch[23].l_um_iw[236] ,
    \top_I.branch[23].l_um_iw[235] ,
    \top_I.branch[23].l_um_iw[234] ,
    \top_I.branch[23].l_um_iw[233] ,
    \top_I.branch[23].l_um_iw[232] ,
    \top_I.branch[23].l_um_iw[231] ,
    \top_I.branch[23].l_um_iw[230] ,
    \top_I.branch[23].l_um_iw[229] ,
    \top_I.branch[23].l_um_iw[228] ,
    \top_I.branch[23].l_um_iw[227] ,
    \top_I.branch[23].l_um_iw[226] ,
    \top_I.branch[23].l_um_iw[225] ,
    \top_I.branch[23].l_um_iw[224] ,
    \top_I.branch[23].l_um_iw[223] ,
    \top_I.branch[23].l_um_iw[222] ,
    \top_I.branch[23].l_um_iw[221] ,
    \top_I.branch[23].l_um_iw[220] ,
    \top_I.branch[23].l_um_iw[219] ,
    \top_I.branch[23].l_um_iw[218] ,
    \top_I.branch[23].l_um_iw[217] ,
    \top_I.branch[23].l_um_iw[216] ,
    \top_I.branch[23].l_um_iw[215] ,
    \top_I.branch[23].l_um_iw[214] ,
    \top_I.branch[23].l_um_iw[213] ,
    \top_I.branch[23].l_um_iw[212] ,
    \top_I.branch[23].l_um_iw[211] ,
    \top_I.branch[23].l_um_iw[210] ,
    \top_I.branch[23].l_um_iw[209] ,
    \top_I.branch[23].l_um_iw[208] ,
    \top_I.branch[23].l_um_iw[207] ,
    \top_I.branch[23].l_um_iw[206] ,
    \top_I.branch[23].l_um_iw[205] ,
    \top_I.branch[23].l_um_iw[204] ,
    \top_I.branch[23].l_um_iw[203] ,
    \top_I.branch[23].l_um_iw[202] ,
    \top_I.branch[23].l_um_iw[201] ,
    \top_I.branch[23].l_um_iw[200] ,
    \top_I.branch[23].l_um_iw[199] ,
    \top_I.branch[23].l_um_iw[198] ,
    \top_I.branch[23].l_um_iw[197] ,
    \top_I.branch[23].l_um_iw[196] ,
    \top_I.branch[23].l_um_iw[195] ,
    \top_I.branch[23].l_um_iw[194] ,
    \top_I.branch[23].l_um_iw[193] ,
    \top_I.branch[23].l_um_iw[192] ,
    \top_I.branch[23].l_um_iw[191] ,
    \top_I.branch[23].l_um_iw[190] ,
    \top_I.branch[23].l_um_iw[189] ,
    \top_I.branch[23].l_um_iw[188] ,
    \top_I.branch[23].l_um_iw[187] ,
    \top_I.branch[23].l_um_iw[186] ,
    \top_I.branch[23].l_um_iw[185] ,
    \top_I.branch[23].l_um_iw[184] ,
    \top_I.branch[23].l_um_iw[183] ,
    \top_I.branch[23].l_um_iw[182] ,
    \top_I.branch[23].l_um_iw[181] ,
    \top_I.branch[23].l_um_iw[180] ,
    \top_I.branch[23].l_um_iw[179] ,
    \top_I.branch[23].l_um_iw[178] ,
    \top_I.branch[23].l_um_iw[177] ,
    \top_I.branch[23].l_um_iw[176] ,
    \top_I.branch[23].l_um_iw[175] ,
    \top_I.branch[23].l_um_iw[174] ,
    \top_I.branch[23].l_um_iw[173] ,
    \top_I.branch[23].l_um_iw[172] ,
    \top_I.branch[23].l_um_iw[171] ,
    \top_I.branch[23].l_um_iw[170] ,
    \top_I.branch[23].l_um_iw[169] ,
    \top_I.branch[23].l_um_iw[168] ,
    \top_I.branch[23].l_um_iw[167] ,
    \top_I.branch[23].l_um_iw[166] ,
    \top_I.branch[23].l_um_iw[165] ,
    \top_I.branch[23].l_um_iw[164] ,
    \top_I.branch[23].l_um_iw[163] ,
    \top_I.branch[23].l_um_iw[162] ,
    \top_I.branch[23].l_um_iw[161] ,
    \top_I.branch[23].l_um_iw[160] ,
    \top_I.branch[23].l_um_iw[159] ,
    \top_I.branch[23].l_um_iw[158] ,
    \top_I.branch[23].l_um_iw[157] ,
    \top_I.branch[23].l_um_iw[156] ,
    \top_I.branch[23].l_um_iw[155] ,
    \top_I.branch[23].l_um_iw[154] ,
    \top_I.branch[23].l_um_iw[153] ,
    \top_I.branch[23].l_um_iw[152] ,
    \top_I.branch[23].l_um_iw[151] ,
    \top_I.branch[23].l_um_iw[150] ,
    \top_I.branch[23].l_um_iw[149] ,
    \top_I.branch[23].l_um_iw[148] ,
    \top_I.branch[23].l_um_iw[147] ,
    \top_I.branch[23].l_um_iw[146] ,
    \top_I.branch[23].l_um_iw[145] ,
    \top_I.branch[23].l_um_iw[144] ,
    \top_I.branch[23].l_um_iw[143] ,
    \top_I.branch[23].l_um_iw[142] ,
    \top_I.branch[23].l_um_iw[141] ,
    \top_I.branch[23].l_um_iw[140] ,
    \top_I.branch[23].l_um_iw[139] ,
    \top_I.branch[23].l_um_iw[138] ,
    \top_I.branch[23].l_um_iw[137] ,
    \top_I.branch[23].l_um_iw[136] ,
    \top_I.branch[23].l_um_iw[135] ,
    \top_I.branch[23].l_um_iw[134] ,
    \top_I.branch[23].l_um_iw[133] ,
    \top_I.branch[23].l_um_iw[132] ,
    \top_I.branch[23].l_um_iw[131] ,
    \top_I.branch[23].l_um_iw[130] ,
    \top_I.branch[23].l_um_iw[129] ,
    \top_I.branch[23].l_um_iw[128] ,
    \top_I.branch[23].l_um_iw[127] ,
    \top_I.branch[23].l_um_iw[126] ,
    \top_I.branch[23].l_um_iw[125] ,
    \top_I.branch[23].l_um_iw[124] ,
    \top_I.branch[23].l_um_iw[123] ,
    \top_I.branch[23].l_um_iw[122] ,
    \top_I.branch[23].l_um_iw[121] ,
    \top_I.branch[23].l_um_iw[120] ,
    \top_I.branch[23].l_um_iw[119] ,
    \top_I.branch[23].l_um_iw[118] ,
    \top_I.branch[23].l_um_iw[117] ,
    \top_I.branch[23].l_um_iw[116] ,
    \top_I.branch[23].l_um_iw[115] ,
    \top_I.branch[23].l_um_iw[114] ,
    \top_I.branch[23].l_um_iw[113] ,
    \top_I.branch[23].l_um_iw[112] ,
    \top_I.branch[23].l_um_iw[111] ,
    \top_I.branch[23].l_um_iw[110] ,
    \top_I.branch[23].l_um_iw[109] ,
    \top_I.branch[23].l_um_iw[108] ,
    \top_I.branch[23].l_um_iw[107] ,
    \top_I.branch[23].l_um_iw[106] ,
    \top_I.branch[23].l_um_iw[105] ,
    \top_I.branch[23].l_um_iw[104] ,
    \top_I.branch[23].l_um_iw[103] ,
    \top_I.branch[23].l_um_iw[102] ,
    \top_I.branch[23].l_um_iw[101] ,
    \top_I.branch[23].l_um_iw[100] ,
    \top_I.branch[23].l_um_iw[99] ,
    \top_I.branch[23].l_um_iw[98] ,
    \top_I.branch[23].l_um_iw[97] ,
    \top_I.branch[23].l_um_iw[96] ,
    \top_I.branch[23].l_um_iw[95] ,
    \top_I.branch[23].l_um_iw[94] ,
    \top_I.branch[23].l_um_iw[93] ,
    \top_I.branch[23].l_um_iw[92] ,
    \top_I.branch[23].l_um_iw[91] ,
    \top_I.branch[23].l_um_iw[90] ,
    \top_I.branch[23].l_um_iw[89] ,
    \top_I.branch[23].l_um_iw[88] ,
    \top_I.branch[23].l_um_iw[87] ,
    \top_I.branch[23].l_um_iw[86] ,
    \top_I.branch[23].l_um_iw[85] ,
    \top_I.branch[23].l_um_iw[84] ,
    \top_I.branch[23].l_um_iw[83] ,
    \top_I.branch[23].l_um_iw[82] ,
    \top_I.branch[23].l_um_iw[81] ,
    \top_I.branch[23].l_um_iw[80] ,
    \top_I.branch[23].l_um_iw[79] ,
    \top_I.branch[23].l_um_iw[78] ,
    \top_I.branch[23].l_um_iw[77] ,
    \top_I.branch[23].l_um_iw[76] ,
    \top_I.branch[23].l_um_iw[75] ,
    \top_I.branch[23].l_um_iw[74] ,
    \top_I.branch[23].l_um_iw[73] ,
    \top_I.branch[23].l_um_iw[72] ,
    \top_I.branch[23].l_um_iw[71] ,
    \top_I.branch[23].l_um_iw[70] ,
    \top_I.branch[23].l_um_iw[69] ,
    \top_I.branch[23].l_um_iw[68] ,
    \top_I.branch[23].l_um_iw[67] ,
    \top_I.branch[23].l_um_iw[66] ,
    \top_I.branch[23].l_um_iw[65] ,
    \top_I.branch[23].l_um_iw[64] ,
    \top_I.branch[23].l_um_iw[63] ,
    \top_I.branch[23].l_um_iw[62] ,
    \top_I.branch[23].l_um_iw[61] ,
    \top_I.branch[23].l_um_iw[60] ,
    \top_I.branch[23].l_um_iw[59] ,
    \top_I.branch[23].l_um_iw[58] ,
    \top_I.branch[23].l_um_iw[57] ,
    \top_I.branch[23].l_um_iw[56] ,
    \top_I.branch[23].l_um_iw[55] ,
    \top_I.branch[23].l_um_iw[54] ,
    \top_I.branch[23].l_um_iw[53] ,
    \top_I.branch[23].l_um_iw[52] ,
    \top_I.branch[23].l_um_iw[51] ,
    \top_I.branch[23].l_um_iw[50] ,
    \top_I.branch[23].l_um_iw[49] ,
    \top_I.branch[23].l_um_iw[48] ,
    \top_I.branch[23].l_um_iw[47] ,
    \top_I.branch[23].l_um_iw[46] ,
    \top_I.branch[23].l_um_iw[45] ,
    \top_I.branch[23].l_um_iw[44] ,
    \top_I.branch[23].l_um_iw[43] ,
    \top_I.branch[23].l_um_iw[42] ,
    \top_I.branch[23].l_um_iw[41] ,
    \top_I.branch[23].l_um_iw[40] ,
    \top_I.branch[23].l_um_iw[39] ,
    \top_I.branch[23].l_um_iw[38] ,
    \top_I.branch[23].l_um_iw[37] ,
    \top_I.branch[23].l_um_iw[36] ,
    \top_I.branch[23].l_um_iw[35] ,
    \top_I.branch[23].l_um_iw[34] ,
    \top_I.branch[23].l_um_iw[33] ,
    \top_I.branch[23].l_um_iw[32] ,
    \top_I.branch[23].l_um_iw[31] ,
    \top_I.branch[23].l_um_iw[30] ,
    \top_I.branch[23].l_um_iw[29] ,
    \top_I.branch[23].l_um_iw[28] ,
    \top_I.branch[23].l_um_iw[27] ,
    \top_I.branch[23].l_um_iw[26] ,
    \top_I.branch[23].l_um_iw[25] ,
    \top_I.branch[23].l_um_iw[24] ,
    \top_I.branch[23].l_um_iw[23] ,
    \top_I.branch[23].l_um_iw[22] ,
    \top_I.branch[23].l_um_iw[21] ,
    \top_I.branch[23].l_um_iw[20] ,
    \top_I.branch[23].l_um_iw[19] ,
    \top_I.branch[23].l_um_iw[18] ,
    \top_I.branch[23].l_um_iw[17] ,
    \top_I.branch[23].l_um_iw[16] ,
    \top_I.branch[23].l_um_iw[15] ,
    \top_I.branch[23].l_um_iw[14] ,
    \top_I.branch[23].l_um_iw[13] ,
    \top_I.branch[23].l_um_iw[12] ,
    \top_I.branch[23].l_um_iw[11] ,
    \top_I.branch[23].l_um_iw[10] ,
    \top_I.branch[23].l_um_iw[9] ,
    \top_I.branch[23].l_um_iw[8] ,
    \top_I.branch[23].l_um_iw[7] ,
    \top_I.branch[23].l_um_iw[6] ,
    \top_I.branch[23].l_um_iw[5] ,
    \top_I.branch[23].l_um_iw[4] ,
    \top_I.branch[23].l_um_iw[3] ,
    \top_I.branch[23].l_um_iw[2] ,
    \top_I.branch[23].l_um_iw[1] ,
    \top_I.branch[23].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[1] ,
    \top_I.branch[23].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[15] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[14] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[13] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[12] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[11] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[10] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[9] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[8] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[7] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[6] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[5] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[4] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[3] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].l_um_k_zero[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[23].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] ,
    \top_I.branch[23].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[2].col_um[0].um_top_I.block_3_0.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[18] ),
    .ena(\top_I.branch[2].l_um_ena[1] ),
    .rst_n(\top_I.branch[2].l_um_iw[19] ),
    .ui_in({\top_I.branch[2].l_um_iw[27] ,
    \top_I.branch[2].l_um_iw[26] ,
    \top_I.branch[2].l_um_iw[25] ,
    \top_I.branch[2].l_um_iw[24] ,
    \top_I.branch[2].l_um_iw[23] ,
    \top_I.branch[2].l_um_iw[22] ,
    \top_I.branch[2].l_um_iw[21] ,
    \top_I.branch[2].l_um_iw[20] }),
    .uio_in({\top_I.branch[2].l_um_iw[35] ,
    \top_I.branch[2].l_um_iw[34] ,
    \top_I.branch[2].l_um_iw[33] ,
    \top_I.branch[2].l_um_iw[32] ,
    \top_I.branch[2].l_um_iw[31] ,
    \top_I.branch[2].l_um_iw[30] ,
    \top_I.branch[2].l_um_iw[29] ,
    \top_I.branch[2].l_um_iw[28] }),
    .uio_oe({\top_I.branch[2].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[0] }));
 tt_um_vga_clock \top_I.branch[2].col_um[1].um_top_I.block_3_1.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[54] ),
    .ena(\top_I.branch[2].l_um_ena[3] ),
    .rst_n(\top_I.branch[2].l_um_iw[55] ),
    .ui_in({\top_I.branch[2].l_um_iw[63] ,
    \top_I.branch[2].l_um_iw[62] ,
    \top_I.branch[2].l_um_iw[61] ,
    \top_I.branch[2].l_um_iw[60] ,
    \top_I.branch[2].l_um_iw[59] ,
    \top_I.branch[2].l_um_iw[58] ,
    \top_I.branch[2].l_um_iw[57] ,
    \top_I.branch[2].l_um_iw[56] }),
    .uio_in({\top_I.branch[2].l_um_iw[71] ,
    \top_I.branch[2].l_um_iw[70] ,
    \top_I.branch[2].l_um_iw[69] ,
    \top_I.branch[2].l_um_iw[68] ,
    \top_I.branch[2].l_um_iw[67] ,
    \top_I.branch[2].l_um_iw[66] ,
    \top_I.branch[2].l_um_iw[65] ,
    \top_I.branch[2].l_um_iw[64] }),
    .uio_oe({\top_I.branch[2].col_um[1].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[1].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[1].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[0] }));
 tt_um_MichaelBell_hovalaag \top_I.branch[2].col_um[2].um_top_I.block_3_2.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[90] ),
    .ena(\top_I.branch[2].l_um_ena[5] ),
    .rst_n(\top_I.branch[2].l_um_iw[91] ),
    .ui_in({\top_I.branch[2].l_um_iw[99] ,
    \top_I.branch[2].l_um_iw[98] ,
    \top_I.branch[2].l_um_iw[97] ,
    \top_I.branch[2].l_um_iw[96] ,
    \top_I.branch[2].l_um_iw[95] ,
    \top_I.branch[2].l_um_iw[94] ,
    \top_I.branch[2].l_um_iw[93] ,
    \top_I.branch[2].l_um_iw[92] }),
    .uio_in({\top_I.branch[2].l_um_iw[107] ,
    \top_I.branch[2].l_um_iw[106] ,
    \top_I.branch[2].l_um_iw[105] ,
    \top_I.branch[2].l_um_iw[104] ,
    \top_I.branch[2].l_um_iw[103] ,
    \top_I.branch[2].l_um_iw[102] ,
    \top_I.branch[2].l_um_iw[101] ,
    \top_I.branch[2].l_um_iw[100] }),
    .uio_oe({\top_I.branch[2].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[0] }));
 tt_um_gatecat_fpga_top \top_I.branch[2].col_um[3].um_top_I.block_3_3.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[126] ),
    .ena(\top_I.branch[2].l_um_ena[7] ),
    .rst_n(\top_I.branch[2].l_um_iw[127] ),
    .ui_in({\top_I.branch[2].l_um_iw[135] ,
    \top_I.branch[2].l_um_iw[134] ,
    \top_I.branch[2].l_um_iw[133] ,
    \top_I.branch[2].l_um_iw[132] ,
    \top_I.branch[2].l_um_iw[131] ,
    \top_I.branch[2].l_um_iw[130] ,
    \top_I.branch[2].l_um_iw[129] ,
    \top_I.branch[2].l_um_iw[128] }),
    .uio_in({\top_I.branch[2].l_um_iw[143] ,
    \top_I.branch[2].l_um_iw[142] ,
    \top_I.branch[2].l_um_iw[141] ,
    \top_I.branch[2].l_um_iw[140] ,
    \top_I.branch[2].l_um_iw[139] ,
    \top_I.branch[2].l_um_iw[138] ,
    \top_I.branch[2].l_um_iw[137] ,
    \top_I.branch[2].l_um_iw[136] }),
    .uio_oe({\top_I.branch[2].col_um[3].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[3].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[3].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[0] }));
 tt_um_millerresearch_top \top_I.branch[2].col_um[4].um_top_I.block_3_4.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[162] ),
    .ena(\top_I.branch[2].l_um_ena[9] ),
    .rst_n(\top_I.branch[2].l_um_iw[163] ),
    .ui_in({\top_I.branch[2].l_um_iw[171] ,
    \top_I.branch[2].l_um_iw[170] ,
    \top_I.branch[2].l_um_iw[169] ,
    \top_I.branch[2].l_um_iw[168] ,
    \top_I.branch[2].l_um_iw[167] ,
    \top_I.branch[2].l_um_iw[166] ,
    \top_I.branch[2].l_um_iw[165] ,
    \top_I.branch[2].l_um_iw[164] }),
    .uio_in({\top_I.branch[2].l_um_iw[179] ,
    \top_I.branch[2].l_um_iw[178] ,
    \top_I.branch[2].l_um_iw[177] ,
    \top_I.branch[2].l_um_iw[176] ,
    \top_I.branch[2].l_um_iw[175] ,
    \top_I.branch[2].l_um_iw[174] ,
    \top_I.branch[2].l_um_iw[173] ,
    \top_I.branch[2].l_um_iw[172] }),
    .uio_oe({\top_I.branch[2].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[0] }));
 tt_um_ringosc_cnt \top_I.branch[2].col_um[5].um_top_I.block_3_5.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[198] ),
    .ena(\top_I.branch[2].l_um_ena[11] ),
    .rst_n(\top_I.branch[2].l_um_iw[199] ),
    .ui_in({\top_I.branch[2].l_um_iw[207] ,
    \top_I.branch[2].l_um_iw[206] ,
    \top_I.branch[2].l_um_iw[205] ,
    \top_I.branch[2].l_um_iw[204] ,
    \top_I.branch[2].l_um_iw[203] ,
    \top_I.branch[2].l_um_iw[202] ,
    \top_I.branch[2].l_um_iw[201] ,
    \top_I.branch[2].l_um_iw[200] }),
    .uio_in({\top_I.branch[2].l_um_iw[215] ,
    \top_I.branch[2].l_um_iw[214] ,
    \top_I.branch[2].l_um_iw[213] ,
    \top_I.branch[2].l_um_iw[212] ,
    \top_I.branch[2].l_um_iw[211] ,
    \top_I.branch[2].l_um_iw[210] ,
    \top_I.branch[2].l_um_iw[209] ,
    \top_I.branch[2].l_um_iw[208] }),
    .uio_oe({\top_I.branch[2].col_um[5].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[5].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[5].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[0] }));
 tt_um_test \top_I.branch[2].col_um[6].um_top_I.block_3_6.tt_um_I  (.clk(\top_I.branch[2].l_um_iw[234] ),
    .ena(\top_I.branch[2].l_um_ena[13] ),
    .rst_n(\top_I.branch[2].l_um_iw[235] ),
    .ui_in({\top_I.branch[2].l_um_iw[243] ,
    \top_I.branch[2].l_um_iw[242] ,
    \top_I.branch[2].l_um_iw[241] ,
    \top_I.branch[2].l_um_iw[240] ,
    \top_I.branch[2].l_um_iw[239] ,
    \top_I.branch[2].l_um_iw[238] ,
    \top_I.branch[2].l_um_iw[237] ,
    \top_I.branch[2].l_um_iw[236] }),
    .uio_in({\top_I.branch[2].l_um_iw[251] ,
    \top_I.branch[2].l_um_iw[250] ,
    \top_I.branch[2].l_um_iw[249] ,
    \top_I.branch[2].l_um_iw[248] ,
    \top_I.branch[2].l_um_iw[247] ,
    \top_I.branch[2].l_um_iw[246] ,
    \top_I.branch[2].l_um_iw[245] ,
    \top_I.branch[2].l_um_iw[244] }),
    .uio_oe({\top_I.branch[2].col_um[6].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[2].col_um[6].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[2].col_um[6].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[2].mux_I  (.k_one(\top_I.branch[2].l_k_one ),
    .k_zero(\top_I.branch[2].l_k_zero ),
    .addr({\top_I.branch[2].l_k_zero ,
    \top_I.branch[2].l_k_zero ,
    \top_I.branch[2].l_k_zero ,
    \top_I.branch[2].l_k_one ,
    \top_I.branch[2].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[2].l_um_ena[15] ,
    \top_I.branch[2].l_um_ena[14] ,
    \top_I.branch[2].l_um_ena[13] ,
    \top_I.branch[2].l_um_ena[12] ,
    \top_I.branch[2].l_um_ena[11] ,
    \top_I.branch[2].l_um_ena[10] ,
    \top_I.branch[2].l_um_ena[9] ,
    \top_I.branch[2].l_um_ena[8] ,
    \top_I.branch[2].l_um_ena[7] ,
    \top_I.branch[2].l_um_ena[6] ,
    \top_I.branch[2].l_um_ena[5] ,
    \top_I.branch[2].l_um_ena[4] ,
    \top_I.branch[2].l_um_ena[3] ,
    \top_I.branch[2].l_um_ena[2] ,
    \top_I.branch[2].l_um_ena[1] ,
    \top_I.branch[2].l_um_ena[0] }),
    .um_iw({\top_I.branch[2].l_um_iw[287] ,
    \top_I.branch[2].l_um_iw[286] ,
    \top_I.branch[2].l_um_iw[285] ,
    \top_I.branch[2].l_um_iw[284] ,
    \top_I.branch[2].l_um_iw[283] ,
    \top_I.branch[2].l_um_iw[282] ,
    \top_I.branch[2].l_um_iw[281] ,
    \top_I.branch[2].l_um_iw[280] ,
    \top_I.branch[2].l_um_iw[279] ,
    \top_I.branch[2].l_um_iw[278] ,
    \top_I.branch[2].l_um_iw[277] ,
    \top_I.branch[2].l_um_iw[276] ,
    \top_I.branch[2].l_um_iw[275] ,
    \top_I.branch[2].l_um_iw[274] ,
    \top_I.branch[2].l_um_iw[273] ,
    \top_I.branch[2].l_um_iw[272] ,
    \top_I.branch[2].l_um_iw[271] ,
    \top_I.branch[2].l_um_iw[270] ,
    \top_I.branch[2].l_um_iw[269] ,
    \top_I.branch[2].l_um_iw[268] ,
    \top_I.branch[2].l_um_iw[267] ,
    \top_I.branch[2].l_um_iw[266] ,
    \top_I.branch[2].l_um_iw[265] ,
    \top_I.branch[2].l_um_iw[264] ,
    \top_I.branch[2].l_um_iw[263] ,
    \top_I.branch[2].l_um_iw[262] ,
    \top_I.branch[2].l_um_iw[261] ,
    \top_I.branch[2].l_um_iw[260] ,
    \top_I.branch[2].l_um_iw[259] ,
    \top_I.branch[2].l_um_iw[258] ,
    \top_I.branch[2].l_um_iw[257] ,
    \top_I.branch[2].l_um_iw[256] ,
    \top_I.branch[2].l_um_iw[255] ,
    \top_I.branch[2].l_um_iw[254] ,
    \top_I.branch[2].l_um_iw[253] ,
    \top_I.branch[2].l_um_iw[252] ,
    \top_I.branch[2].l_um_iw[251] ,
    \top_I.branch[2].l_um_iw[250] ,
    \top_I.branch[2].l_um_iw[249] ,
    \top_I.branch[2].l_um_iw[248] ,
    \top_I.branch[2].l_um_iw[247] ,
    \top_I.branch[2].l_um_iw[246] ,
    \top_I.branch[2].l_um_iw[245] ,
    \top_I.branch[2].l_um_iw[244] ,
    \top_I.branch[2].l_um_iw[243] ,
    \top_I.branch[2].l_um_iw[242] ,
    \top_I.branch[2].l_um_iw[241] ,
    \top_I.branch[2].l_um_iw[240] ,
    \top_I.branch[2].l_um_iw[239] ,
    \top_I.branch[2].l_um_iw[238] ,
    \top_I.branch[2].l_um_iw[237] ,
    \top_I.branch[2].l_um_iw[236] ,
    \top_I.branch[2].l_um_iw[235] ,
    \top_I.branch[2].l_um_iw[234] ,
    \top_I.branch[2].l_um_iw[233] ,
    \top_I.branch[2].l_um_iw[232] ,
    \top_I.branch[2].l_um_iw[231] ,
    \top_I.branch[2].l_um_iw[230] ,
    \top_I.branch[2].l_um_iw[229] ,
    \top_I.branch[2].l_um_iw[228] ,
    \top_I.branch[2].l_um_iw[227] ,
    \top_I.branch[2].l_um_iw[226] ,
    \top_I.branch[2].l_um_iw[225] ,
    \top_I.branch[2].l_um_iw[224] ,
    \top_I.branch[2].l_um_iw[223] ,
    \top_I.branch[2].l_um_iw[222] ,
    \top_I.branch[2].l_um_iw[221] ,
    \top_I.branch[2].l_um_iw[220] ,
    \top_I.branch[2].l_um_iw[219] ,
    \top_I.branch[2].l_um_iw[218] ,
    \top_I.branch[2].l_um_iw[217] ,
    \top_I.branch[2].l_um_iw[216] ,
    \top_I.branch[2].l_um_iw[215] ,
    \top_I.branch[2].l_um_iw[214] ,
    \top_I.branch[2].l_um_iw[213] ,
    \top_I.branch[2].l_um_iw[212] ,
    \top_I.branch[2].l_um_iw[211] ,
    \top_I.branch[2].l_um_iw[210] ,
    \top_I.branch[2].l_um_iw[209] ,
    \top_I.branch[2].l_um_iw[208] ,
    \top_I.branch[2].l_um_iw[207] ,
    \top_I.branch[2].l_um_iw[206] ,
    \top_I.branch[2].l_um_iw[205] ,
    \top_I.branch[2].l_um_iw[204] ,
    \top_I.branch[2].l_um_iw[203] ,
    \top_I.branch[2].l_um_iw[202] ,
    \top_I.branch[2].l_um_iw[201] ,
    \top_I.branch[2].l_um_iw[200] ,
    \top_I.branch[2].l_um_iw[199] ,
    \top_I.branch[2].l_um_iw[198] ,
    \top_I.branch[2].l_um_iw[197] ,
    \top_I.branch[2].l_um_iw[196] ,
    \top_I.branch[2].l_um_iw[195] ,
    \top_I.branch[2].l_um_iw[194] ,
    \top_I.branch[2].l_um_iw[193] ,
    \top_I.branch[2].l_um_iw[192] ,
    \top_I.branch[2].l_um_iw[191] ,
    \top_I.branch[2].l_um_iw[190] ,
    \top_I.branch[2].l_um_iw[189] ,
    \top_I.branch[2].l_um_iw[188] ,
    \top_I.branch[2].l_um_iw[187] ,
    \top_I.branch[2].l_um_iw[186] ,
    \top_I.branch[2].l_um_iw[185] ,
    \top_I.branch[2].l_um_iw[184] ,
    \top_I.branch[2].l_um_iw[183] ,
    \top_I.branch[2].l_um_iw[182] ,
    \top_I.branch[2].l_um_iw[181] ,
    \top_I.branch[2].l_um_iw[180] ,
    \top_I.branch[2].l_um_iw[179] ,
    \top_I.branch[2].l_um_iw[178] ,
    \top_I.branch[2].l_um_iw[177] ,
    \top_I.branch[2].l_um_iw[176] ,
    \top_I.branch[2].l_um_iw[175] ,
    \top_I.branch[2].l_um_iw[174] ,
    \top_I.branch[2].l_um_iw[173] ,
    \top_I.branch[2].l_um_iw[172] ,
    \top_I.branch[2].l_um_iw[171] ,
    \top_I.branch[2].l_um_iw[170] ,
    \top_I.branch[2].l_um_iw[169] ,
    \top_I.branch[2].l_um_iw[168] ,
    \top_I.branch[2].l_um_iw[167] ,
    \top_I.branch[2].l_um_iw[166] ,
    \top_I.branch[2].l_um_iw[165] ,
    \top_I.branch[2].l_um_iw[164] ,
    \top_I.branch[2].l_um_iw[163] ,
    \top_I.branch[2].l_um_iw[162] ,
    \top_I.branch[2].l_um_iw[161] ,
    \top_I.branch[2].l_um_iw[160] ,
    \top_I.branch[2].l_um_iw[159] ,
    \top_I.branch[2].l_um_iw[158] ,
    \top_I.branch[2].l_um_iw[157] ,
    \top_I.branch[2].l_um_iw[156] ,
    \top_I.branch[2].l_um_iw[155] ,
    \top_I.branch[2].l_um_iw[154] ,
    \top_I.branch[2].l_um_iw[153] ,
    \top_I.branch[2].l_um_iw[152] ,
    \top_I.branch[2].l_um_iw[151] ,
    \top_I.branch[2].l_um_iw[150] ,
    \top_I.branch[2].l_um_iw[149] ,
    \top_I.branch[2].l_um_iw[148] ,
    \top_I.branch[2].l_um_iw[147] ,
    \top_I.branch[2].l_um_iw[146] ,
    \top_I.branch[2].l_um_iw[145] ,
    \top_I.branch[2].l_um_iw[144] ,
    \top_I.branch[2].l_um_iw[143] ,
    \top_I.branch[2].l_um_iw[142] ,
    \top_I.branch[2].l_um_iw[141] ,
    \top_I.branch[2].l_um_iw[140] ,
    \top_I.branch[2].l_um_iw[139] ,
    \top_I.branch[2].l_um_iw[138] ,
    \top_I.branch[2].l_um_iw[137] ,
    \top_I.branch[2].l_um_iw[136] ,
    \top_I.branch[2].l_um_iw[135] ,
    \top_I.branch[2].l_um_iw[134] ,
    \top_I.branch[2].l_um_iw[133] ,
    \top_I.branch[2].l_um_iw[132] ,
    \top_I.branch[2].l_um_iw[131] ,
    \top_I.branch[2].l_um_iw[130] ,
    \top_I.branch[2].l_um_iw[129] ,
    \top_I.branch[2].l_um_iw[128] ,
    \top_I.branch[2].l_um_iw[127] ,
    \top_I.branch[2].l_um_iw[126] ,
    \top_I.branch[2].l_um_iw[125] ,
    \top_I.branch[2].l_um_iw[124] ,
    \top_I.branch[2].l_um_iw[123] ,
    \top_I.branch[2].l_um_iw[122] ,
    \top_I.branch[2].l_um_iw[121] ,
    \top_I.branch[2].l_um_iw[120] ,
    \top_I.branch[2].l_um_iw[119] ,
    \top_I.branch[2].l_um_iw[118] ,
    \top_I.branch[2].l_um_iw[117] ,
    \top_I.branch[2].l_um_iw[116] ,
    \top_I.branch[2].l_um_iw[115] ,
    \top_I.branch[2].l_um_iw[114] ,
    \top_I.branch[2].l_um_iw[113] ,
    \top_I.branch[2].l_um_iw[112] ,
    \top_I.branch[2].l_um_iw[111] ,
    \top_I.branch[2].l_um_iw[110] ,
    \top_I.branch[2].l_um_iw[109] ,
    \top_I.branch[2].l_um_iw[108] ,
    \top_I.branch[2].l_um_iw[107] ,
    \top_I.branch[2].l_um_iw[106] ,
    \top_I.branch[2].l_um_iw[105] ,
    \top_I.branch[2].l_um_iw[104] ,
    \top_I.branch[2].l_um_iw[103] ,
    \top_I.branch[2].l_um_iw[102] ,
    \top_I.branch[2].l_um_iw[101] ,
    \top_I.branch[2].l_um_iw[100] ,
    \top_I.branch[2].l_um_iw[99] ,
    \top_I.branch[2].l_um_iw[98] ,
    \top_I.branch[2].l_um_iw[97] ,
    \top_I.branch[2].l_um_iw[96] ,
    \top_I.branch[2].l_um_iw[95] ,
    \top_I.branch[2].l_um_iw[94] ,
    \top_I.branch[2].l_um_iw[93] ,
    \top_I.branch[2].l_um_iw[92] ,
    \top_I.branch[2].l_um_iw[91] ,
    \top_I.branch[2].l_um_iw[90] ,
    \top_I.branch[2].l_um_iw[89] ,
    \top_I.branch[2].l_um_iw[88] ,
    \top_I.branch[2].l_um_iw[87] ,
    \top_I.branch[2].l_um_iw[86] ,
    \top_I.branch[2].l_um_iw[85] ,
    \top_I.branch[2].l_um_iw[84] ,
    \top_I.branch[2].l_um_iw[83] ,
    \top_I.branch[2].l_um_iw[82] ,
    \top_I.branch[2].l_um_iw[81] ,
    \top_I.branch[2].l_um_iw[80] ,
    \top_I.branch[2].l_um_iw[79] ,
    \top_I.branch[2].l_um_iw[78] ,
    \top_I.branch[2].l_um_iw[77] ,
    \top_I.branch[2].l_um_iw[76] ,
    \top_I.branch[2].l_um_iw[75] ,
    \top_I.branch[2].l_um_iw[74] ,
    \top_I.branch[2].l_um_iw[73] ,
    \top_I.branch[2].l_um_iw[72] ,
    \top_I.branch[2].l_um_iw[71] ,
    \top_I.branch[2].l_um_iw[70] ,
    \top_I.branch[2].l_um_iw[69] ,
    \top_I.branch[2].l_um_iw[68] ,
    \top_I.branch[2].l_um_iw[67] ,
    \top_I.branch[2].l_um_iw[66] ,
    \top_I.branch[2].l_um_iw[65] ,
    \top_I.branch[2].l_um_iw[64] ,
    \top_I.branch[2].l_um_iw[63] ,
    \top_I.branch[2].l_um_iw[62] ,
    \top_I.branch[2].l_um_iw[61] ,
    \top_I.branch[2].l_um_iw[60] ,
    \top_I.branch[2].l_um_iw[59] ,
    \top_I.branch[2].l_um_iw[58] ,
    \top_I.branch[2].l_um_iw[57] ,
    \top_I.branch[2].l_um_iw[56] ,
    \top_I.branch[2].l_um_iw[55] ,
    \top_I.branch[2].l_um_iw[54] ,
    \top_I.branch[2].l_um_iw[53] ,
    \top_I.branch[2].l_um_iw[52] ,
    \top_I.branch[2].l_um_iw[51] ,
    \top_I.branch[2].l_um_iw[50] ,
    \top_I.branch[2].l_um_iw[49] ,
    \top_I.branch[2].l_um_iw[48] ,
    \top_I.branch[2].l_um_iw[47] ,
    \top_I.branch[2].l_um_iw[46] ,
    \top_I.branch[2].l_um_iw[45] ,
    \top_I.branch[2].l_um_iw[44] ,
    \top_I.branch[2].l_um_iw[43] ,
    \top_I.branch[2].l_um_iw[42] ,
    \top_I.branch[2].l_um_iw[41] ,
    \top_I.branch[2].l_um_iw[40] ,
    \top_I.branch[2].l_um_iw[39] ,
    \top_I.branch[2].l_um_iw[38] ,
    \top_I.branch[2].l_um_iw[37] ,
    \top_I.branch[2].l_um_iw[36] ,
    \top_I.branch[2].l_um_iw[35] ,
    \top_I.branch[2].l_um_iw[34] ,
    \top_I.branch[2].l_um_iw[33] ,
    \top_I.branch[2].l_um_iw[32] ,
    \top_I.branch[2].l_um_iw[31] ,
    \top_I.branch[2].l_um_iw[30] ,
    \top_I.branch[2].l_um_iw[29] ,
    \top_I.branch[2].l_um_iw[28] ,
    \top_I.branch[2].l_um_iw[27] ,
    \top_I.branch[2].l_um_iw[26] ,
    \top_I.branch[2].l_um_iw[25] ,
    \top_I.branch[2].l_um_iw[24] ,
    \top_I.branch[2].l_um_iw[23] ,
    \top_I.branch[2].l_um_iw[22] ,
    \top_I.branch[2].l_um_iw[21] ,
    \top_I.branch[2].l_um_iw[20] ,
    \top_I.branch[2].l_um_iw[19] ,
    \top_I.branch[2].l_um_iw[18] ,
    \top_I.branch[2].l_um_iw[17] ,
    \top_I.branch[2].l_um_iw[16] ,
    \top_I.branch[2].l_um_iw[15] ,
    \top_I.branch[2].l_um_iw[14] ,
    \top_I.branch[2].l_um_iw[13] ,
    \top_I.branch[2].l_um_iw[12] ,
    \top_I.branch[2].l_um_iw[11] ,
    \top_I.branch[2].l_um_iw[10] ,
    \top_I.branch[2].l_um_iw[9] ,
    \top_I.branch[2].l_um_iw[8] ,
    \top_I.branch[2].l_um_iw[7] ,
    \top_I.branch[2].l_um_iw[6] ,
    \top_I.branch[2].l_um_iw[5] ,
    \top_I.branch[2].l_um_iw[4] ,
    \top_I.branch[2].l_um_iw[3] ,
    \top_I.branch[2].l_um_iw[2] ,
    \top_I.branch[2].l_um_iw[1] ,
    \top_I.branch[2].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[13] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[11] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[9] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[7] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[5] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[3] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[1] ,
    \top_I.branch[2].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[15] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].l_um_k_zero[14] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[6].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].l_um_k_zero[12] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[5].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].l_um_k_zero[10] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[4].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].l_um_k_zero[8] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[3].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].l_um_k_zero[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[2].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].l_um_k_zero[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[1].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].l_um_k_zero[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[2].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] ,
    \top_I.branch[2].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[3].col_um[0].um_top_I.block_3_16.tt_um_I  (.clk(\top_I.branch[3].l_um_iw[18] ),
    .ena(\top_I.branch[3].l_um_ena[1] ),
    .rst_n(\top_I.branch[3].l_um_iw[19] ),
    .ui_in({\top_I.branch[3].l_um_iw[27] ,
    \top_I.branch[3].l_um_iw[26] ,
    \top_I.branch[3].l_um_iw[25] ,
    \top_I.branch[3].l_um_iw[24] ,
    \top_I.branch[3].l_um_iw[23] ,
    \top_I.branch[3].l_um_iw[22] ,
    \top_I.branch[3].l_um_iw[21] ,
    \top_I.branch[3].l_um_iw[20] }),
    .uio_in({\top_I.branch[3].l_um_iw[35] ,
    \top_I.branch[3].l_um_iw[34] ,
    \top_I.branch[3].l_um_iw[33] ,
    \top_I.branch[3].l_um_iw[32] ,
    \top_I.branch[3].l_um_iw[31] ,
    \top_I.branch[3].l_um_iw[30] ,
    \top_I.branch[3].l_um_iw[29] ,
    \top_I.branch[3].l_um_iw[28] }),
    .uio_oe({\top_I.branch[3].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[3].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[3].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[3].mux_I  (.k_one(\top_I.branch[3].l_k_one ),
    .k_zero(\top_I.branch[3].l_k_zero ),
    .addr({\top_I.branch[3].l_k_zero ,
    \top_I.branch[3].l_k_zero ,
    \top_I.branch[3].l_k_zero ,
    \top_I.branch[3].l_k_one ,
    \top_I.branch[3].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[3].l_um_ena[15] ,
    \top_I.branch[3].l_um_ena[14] ,
    \top_I.branch[3].l_um_ena[13] ,
    \top_I.branch[3].l_um_ena[12] ,
    \top_I.branch[3].l_um_ena[11] ,
    \top_I.branch[3].l_um_ena[10] ,
    \top_I.branch[3].l_um_ena[9] ,
    \top_I.branch[3].l_um_ena[8] ,
    \top_I.branch[3].l_um_ena[7] ,
    \top_I.branch[3].l_um_ena[6] ,
    \top_I.branch[3].l_um_ena[5] ,
    \top_I.branch[3].l_um_ena[4] ,
    \top_I.branch[3].l_um_ena[3] ,
    \top_I.branch[3].l_um_ena[2] ,
    \top_I.branch[3].l_um_ena[1] ,
    \top_I.branch[3].l_um_ena[0] }),
    .um_iw({\top_I.branch[3].l_um_iw[287] ,
    \top_I.branch[3].l_um_iw[286] ,
    \top_I.branch[3].l_um_iw[285] ,
    \top_I.branch[3].l_um_iw[284] ,
    \top_I.branch[3].l_um_iw[283] ,
    \top_I.branch[3].l_um_iw[282] ,
    \top_I.branch[3].l_um_iw[281] ,
    \top_I.branch[3].l_um_iw[280] ,
    \top_I.branch[3].l_um_iw[279] ,
    \top_I.branch[3].l_um_iw[278] ,
    \top_I.branch[3].l_um_iw[277] ,
    \top_I.branch[3].l_um_iw[276] ,
    \top_I.branch[3].l_um_iw[275] ,
    \top_I.branch[3].l_um_iw[274] ,
    \top_I.branch[3].l_um_iw[273] ,
    \top_I.branch[3].l_um_iw[272] ,
    \top_I.branch[3].l_um_iw[271] ,
    \top_I.branch[3].l_um_iw[270] ,
    \top_I.branch[3].l_um_iw[269] ,
    \top_I.branch[3].l_um_iw[268] ,
    \top_I.branch[3].l_um_iw[267] ,
    \top_I.branch[3].l_um_iw[266] ,
    \top_I.branch[3].l_um_iw[265] ,
    \top_I.branch[3].l_um_iw[264] ,
    \top_I.branch[3].l_um_iw[263] ,
    \top_I.branch[3].l_um_iw[262] ,
    \top_I.branch[3].l_um_iw[261] ,
    \top_I.branch[3].l_um_iw[260] ,
    \top_I.branch[3].l_um_iw[259] ,
    \top_I.branch[3].l_um_iw[258] ,
    \top_I.branch[3].l_um_iw[257] ,
    \top_I.branch[3].l_um_iw[256] ,
    \top_I.branch[3].l_um_iw[255] ,
    \top_I.branch[3].l_um_iw[254] ,
    \top_I.branch[3].l_um_iw[253] ,
    \top_I.branch[3].l_um_iw[252] ,
    \top_I.branch[3].l_um_iw[251] ,
    \top_I.branch[3].l_um_iw[250] ,
    \top_I.branch[3].l_um_iw[249] ,
    \top_I.branch[3].l_um_iw[248] ,
    \top_I.branch[3].l_um_iw[247] ,
    \top_I.branch[3].l_um_iw[246] ,
    \top_I.branch[3].l_um_iw[245] ,
    \top_I.branch[3].l_um_iw[244] ,
    \top_I.branch[3].l_um_iw[243] ,
    \top_I.branch[3].l_um_iw[242] ,
    \top_I.branch[3].l_um_iw[241] ,
    \top_I.branch[3].l_um_iw[240] ,
    \top_I.branch[3].l_um_iw[239] ,
    \top_I.branch[3].l_um_iw[238] ,
    \top_I.branch[3].l_um_iw[237] ,
    \top_I.branch[3].l_um_iw[236] ,
    \top_I.branch[3].l_um_iw[235] ,
    \top_I.branch[3].l_um_iw[234] ,
    \top_I.branch[3].l_um_iw[233] ,
    \top_I.branch[3].l_um_iw[232] ,
    \top_I.branch[3].l_um_iw[231] ,
    \top_I.branch[3].l_um_iw[230] ,
    \top_I.branch[3].l_um_iw[229] ,
    \top_I.branch[3].l_um_iw[228] ,
    \top_I.branch[3].l_um_iw[227] ,
    \top_I.branch[3].l_um_iw[226] ,
    \top_I.branch[3].l_um_iw[225] ,
    \top_I.branch[3].l_um_iw[224] ,
    \top_I.branch[3].l_um_iw[223] ,
    \top_I.branch[3].l_um_iw[222] ,
    \top_I.branch[3].l_um_iw[221] ,
    \top_I.branch[3].l_um_iw[220] ,
    \top_I.branch[3].l_um_iw[219] ,
    \top_I.branch[3].l_um_iw[218] ,
    \top_I.branch[3].l_um_iw[217] ,
    \top_I.branch[3].l_um_iw[216] ,
    \top_I.branch[3].l_um_iw[215] ,
    \top_I.branch[3].l_um_iw[214] ,
    \top_I.branch[3].l_um_iw[213] ,
    \top_I.branch[3].l_um_iw[212] ,
    \top_I.branch[3].l_um_iw[211] ,
    \top_I.branch[3].l_um_iw[210] ,
    \top_I.branch[3].l_um_iw[209] ,
    \top_I.branch[3].l_um_iw[208] ,
    \top_I.branch[3].l_um_iw[207] ,
    \top_I.branch[3].l_um_iw[206] ,
    \top_I.branch[3].l_um_iw[205] ,
    \top_I.branch[3].l_um_iw[204] ,
    \top_I.branch[3].l_um_iw[203] ,
    \top_I.branch[3].l_um_iw[202] ,
    \top_I.branch[3].l_um_iw[201] ,
    \top_I.branch[3].l_um_iw[200] ,
    \top_I.branch[3].l_um_iw[199] ,
    \top_I.branch[3].l_um_iw[198] ,
    \top_I.branch[3].l_um_iw[197] ,
    \top_I.branch[3].l_um_iw[196] ,
    \top_I.branch[3].l_um_iw[195] ,
    \top_I.branch[3].l_um_iw[194] ,
    \top_I.branch[3].l_um_iw[193] ,
    \top_I.branch[3].l_um_iw[192] ,
    \top_I.branch[3].l_um_iw[191] ,
    \top_I.branch[3].l_um_iw[190] ,
    \top_I.branch[3].l_um_iw[189] ,
    \top_I.branch[3].l_um_iw[188] ,
    \top_I.branch[3].l_um_iw[187] ,
    \top_I.branch[3].l_um_iw[186] ,
    \top_I.branch[3].l_um_iw[185] ,
    \top_I.branch[3].l_um_iw[184] ,
    \top_I.branch[3].l_um_iw[183] ,
    \top_I.branch[3].l_um_iw[182] ,
    \top_I.branch[3].l_um_iw[181] ,
    \top_I.branch[3].l_um_iw[180] ,
    \top_I.branch[3].l_um_iw[179] ,
    \top_I.branch[3].l_um_iw[178] ,
    \top_I.branch[3].l_um_iw[177] ,
    \top_I.branch[3].l_um_iw[176] ,
    \top_I.branch[3].l_um_iw[175] ,
    \top_I.branch[3].l_um_iw[174] ,
    \top_I.branch[3].l_um_iw[173] ,
    \top_I.branch[3].l_um_iw[172] ,
    \top_I.branch[3].l_um_iw[171] ,
    \top_I.branch[3].l_um_iw[170] ,
    \top_I.branch[3].l_um_iw[169] ,
    \top_I.branch[3].l_um_iw[168] ,
    \top_I.branch[3].l_um_iw[167] ,
    \top_I.branch[3].l_um_iw[166] ,
    \top_I.branch[3].l_um_iw[165] ,
    \top_I.branch[3].l_um_iw[164] ,
    \top_I.branch[3].l_um_iw[163] ,
    \top_I.branch[3].l_um_iw[162] ,
    \top_I.branch[3].l_um_iw[161] ,
    \top_I.branch[3].l_um_iw[160] ,
    \top_I.branch[3].l_um_iw[159] ,
    \top_I.branch[3].l_um_iw[158] ,
    \top_I.branch[3].l_um_iw[157] ,
    \top_I.branch[3].l_um_iw[156] ,
    \top_I.branch[3].l_um_iw[155] ,
    \top_I.branch[3].l_um_iw[154] ,
    \top_I.branch[3].l_um_iw[153] ,
    \top_I.branch[3].l_um_iw[152] ,
    \top_I.branch[3].l_um_iw[151] ,
    \top_I.branch[3].l_um_iw[150] ,
    \top_I.branch[3].l_um_iw[149] ,
    \top_I.branch[3].l_um_iw[148] ,
    \top_I.branch[3].l_um_iw[147] ,
    \top_I.branch[3].l_um_iw[146] ,
    \top_I.branch[3].l_um_iw[145] ,
    \top_I.branch[3].l_um_iw[144] ,
    \top_I.branch[3].l_um_iw[143] ,
    \top_I.branch[3].l_um_iw[142] ,
    \top_I.branch[3].l_um_iw[141] ,
    \top_I.branch[3].l_um_iw[140] ,
    \top_I.branch[3].l_um_iw[139] ,
    \top_I.branch[3].l_um_iw[138] ,
    \top_I.branch[3].l_um_iw[137] ,
    \top_I.branch[3].l_um_iw[136] ,
    \top_I.branch[3].l_um_iw[135] ,
    \top_I.branch[3].l_um_iw[134] ,
    \top_I.branch[3].l_um_iw[133] ,
    \top_I.branch[3].l_um_iw[132] ,
    \top_I.branch[3].l_um_iw[131] ,
    \top_I.branch[3].l_um_iw[130] ,
    \top_I.branch[3].l_um_iw[129] ,
    \top_I.branch[3].l_um_iw[128] ,
    \top_I.branch[3].l_um_iw[127] ,
    \top_I.branch[3].l_um_iw[126] ,
    \top_I.branch[3].l_um_iw[125] ,
    \top_I.branch[3].l_um_iw[124] ,
    \top_I.branch[3].l_um_iw[123] ,
    \top_I.branch[3].l_um_iw[122] ,
    \top_I.branch[3].l_um_iw[121] ,
    \top_I.branch[3].l_um_iw[120] ,
    \top_I.branch[3].l_um_iw[119] ,
    \top_I.branch[3].l_um_iw[118] ,
    \top_I.branch[3].l_um_iw[117] ,
    \top_I.branch[3].l_um_iw[116] ,
    \top_I.branch[3].l_um_iw[115] ,
    \top_I.branch[3].l_um_iw[114] ,
    \top_I.branch[3].l_um_iw[113] ,
    \top_I.branch[3].l_um_iw[112] ,
    \top_I.branch[3].l_um_iw[111] ,
    \top_I.branch[3].l_um_iw[110] ,
    \top_I.branch[3].l_um_iw[109] ,
    \top_I.branch[3].l_um_iw[108] ,
    \top_I.branch[3].l_um_iw[107] ,
    \top_I.branch[3].l_um_iw[106] ,
    \top_I.branch[3].l_um_iw[105] ,
    \top_I.branch[3].l_um_iw[104] ,
    \top_I.branch[3].l_um_iw[103] ,
    \top_I.branch[3].l_um_iw[102] ,
    \top_I.branch[3].l_um_iw[101] ,
    \top_I.branch[3].l_um_iw[100] ,
    \top_I.branch[3].l_um_iw[99] ,
    \top_I.branch[3].l_um_iw[98] ,
    \top_I.branch[3].l_um_iw[97] ,
    \top_I.branch[3].l_um_iw[96] ,
    \top_I.branch[3].l_um_iw[95] ,
    \top_I.branch[3].l_um_iw[94] ,
    \top_I.branch[3].l_um_iw[93] ,
    \top_I.branch[3].l_um_iw[92] ,
    \top_I.branch[3].l_um_iw[91] ,
    \top_I.branch[3].l_um_iw[90] ,
    \top_I.branch[3].l_um_iw[89] ,
    \top_I.branch[3].l_um_iw[88] ,
    \top_I.branch[3].l_um_iw[87] ,
    \top_I.branch[3].l_um_iw[86] ,
    \top_I.branch[3].l_um_iw[85] ,
    \top_I.branch[3].l_um_iw[84] ,
    \top_I.branch[3].l_um_iw[83] ,
    \top_I.branch[3].l_um_iw[82] ,
    \top_I.branch[3].l_um_iw[81] ,
    \top_I.branch[3].l_um_iw[80] ,
    \top_I.branch[3].l_um_iw[79] ,
    \top_I.branch[3].l_um_iw[78] ,
    \top_I.branch[3].l_um_iw[77] ,
    \top_I.branch[3].l_um_iw[76] ,
    \top_I.branch[3].l_um_iw[75] ,
    \top_I.branch[3].l_um_iw[74] ,
    \top_I.branch[3].l_um_iw[73] ,
    \top_I.branch[3].l_um_iw[72] ,
    \top_I.branch[3].l_um_iw[71] ,
    \top_I.branch[3].l_um_iw[70] ,
    \top_I.branch[3].l_um_iw[69] ,
    \top_I.branch[3].l_um_iw[68] ,
    \top_I.branch[3].l_um_iw[67] ,
    \top_I.branch[3].l_um_iw[66] ,
    \top_I.branch[3].l_um_iw[65] ,
    \top_I.branch[3].l_um_iw[64] ,
    \top_I.branch[3].l_um_iw[63] ,
    \top_I.branch[3].l_um_iw[62] ,
    \top_I.branch[3].l_um_iw[61] ,
    \top_I.branch[3].l_um_iw[60] ,
    \top_I.branch[3].l_um_iw[59] ,
    \top_I.branch[3].l_um_iw[58] ,
    \top_I.branch[3].l_um_iw[57] ,
    \top_I.branch[3].l_um_iw[56] ,
    \top_I.branch[3].l_um_iw[55] ,
    \top_I.branch[3].l_um_iw[54] ,
    \top_I.branch[3].l_um_iw[53] ,
    \top_I.branch[3].l_um_iw[52] ,
    \top_I.branch[3].l_um_iw[51] ,
    \top_I.branch[3].l_um_iw[50] ,
    \top_I.branch[3].l_um_iw[49] ,
    \top_I.branch[3].l_um_iw[48] ,
    \top_I.branch[3].l_um_iw[47] ,
    \top_I.branch[3].l_um_iw[46] ,
    \top_I.branch[3].l_um_iw[45] ,
    \top_I.branch[3].l_um_iw[44] ,
    \top_I.branch[3].l_um_iw[43] ,
    \top_I.branch[3].l_um_iw[42] ,
    \top_I.branch[3].l_um_iw[41] ,
    \top_I.branch[3].l_um_iw[40] ,
    \top_I.branch[3].l_um_iw[39] ,
    \top_I.branch[3].l_um_iw[38] ,
    \top_I.branch[3].l_um_iw[37] ,
    \top_I.branch[3].l_um_iw[36] ,
    \top_I.branch[3].l_um_iw[35] ,
    \top_I.branch[3].l_um_iw[34] ,
    \top_I.branch[3].l_um_iw[33] ,
    \top_I.branch[3].l_um_iw[32] ,
    \top_I.branch[3].l_um_iw[31] ,
    \top_I.branch[3].l_um_iw[30] ,
    \top_I.branch[3].l_um_iw[29] ,
    \top_I.branch[3].l_um_iw[28] ,
    \top_I.branch[3].l_um_iw[27] ,
    \top_I.branch[3].l_um_iw[26] ,
    \top_I.branch[3].l_um_iw[25] ,
    \top_I.branch[3].l_um_iw[24] ,
    \top_I.branch[3].l_um_iw[23] ,
    \top_I.branch[3].l_um_iw[22] ,
    \top_I.branch[3].l_um_iw[21] ,
    \top_I.branch[3].l_um_iw[20] ,
    \top_I.branch[3].l_um_iw[19] ,
    \top_I.branch[3].l_um_iw[18] ,
    \top_I.branch[3].l_um_iw[17] ,
    \top_I.branch[3].l_um_iw[16] ,
    \top_I.branch[3].l_um_iw[15] ,
    \top_I.branch[3].l_um_iw[14] ,
    \top_I.branch[3].l_um_iw[13] ,
    \top_I.branch[3].l_um_iw[12] ,
    \top_I.branch[3].l_um_iw[11] ,
    \top_I.branch[3].l_um_iw[10] ,
    \top_I.branch[3].l_um_iw[9] ,
    \top_I.branch[3].l_um_iw[8] ,
    \top_I.branch[3].l_um_iw[7] ,
    \top_I.branch[3].l_um_iw[6] ,
    \top_I.branch[3].l_um_iw[5] ,
    \top_I.branch[3].l_um_iw[4] ,
    \top_I.branch[3].l_um_iw[3] ,
    \top_I.branch[3].l_um_iw[2] ,
    \top_I.branch[3].l_um_iw[1] ,
    \top_I.branch[3].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[1] ,
    \top_I.branch[3].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[15] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[14] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[13] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[12] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[11] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[10] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[9] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[8] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[7] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[6] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[5] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[4] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[3] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].l_um_k_zero[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[3].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] ,
    \top_I.branch[3].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[4].col_um[0].um_bot_I.block_4_0.tt_um_I  (.clk(\top_I.branch[4].l_um_iw[0] ),
    .ena(\top_I.branch[4].l_um_ena[0] ),
    .rst_n(\top_I.branch[4].l_um_iw[1] ),
    .ui_in({\top_I.branch[4].l_um_iw[9] ,
    \top_I.branch[4].l_um_iw[8] ,
    \top_I.branch[4].l_um_iw[7] ,
    \top_I.branch[4].l_um_iw[6] ,
    \top_I.branch[4].l_um_iw[5] ,
    \top_I.branch[4].l_um_iw[4] ,
    \top_I.branch[4].l_um_iw[3] ,
    \top_I.branch[4].l_um_iw[2] }),
    .uio_in({\top_I.branch[4].l_um_iw[17] ,
    \top_I.branch[4].l_um_iw[16] ,
    \top_I.branch[4].l_um_iw[15] ,
    \top_I.branch[4].l_um_iw[14] ,
    \top_I.branch[4].l_um_iw[13] ,
    \top_I.branch[4].l_um_iw[12] ,
    \top_I.branch[4].l_um_iw[11] ,
    \top_I.branch[4].l_um_iw[10] }),
    .uio_oe({\top_I.branch[4].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[4].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[4].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_greycode_top \top_I.branch[4].col_um[2].um_top_I.block_5_2.tt_um_I  (.clk(\top_I.branch[4].l_um_iw[90] ),
    .ena(\top_I.branch[4].l_um_ena[5] ),
    .rst_n(\top_I.branch[4].l_um_iw[91] ),
    .ui_in({\top_I.branch[4].l_um_iw[99] ,
    \top_I.branch[4].l_um_iw[98] ,
    \top_I.branch[4].l_um_iw[97] ,
    \top_I.branch[4].l_um_iw[96] ,
    \top_I.branch[4].l_um_iw[95] ,
    \top_I.branch[4].l_um_iw[94] ,
    \top_I.branch[4].l_um_iw[93] ,
    \top_I.branch[4].l_um_iw[92] }),
    .uio_in({\top_I.branch[4].l_um_iw[107] ,
    \top_I.branch[4].l_um_iw[106] ,
    \top_I.branch[4].l_um_iw[105] ,
    \top_I.branch[4].l_um_iw[104] ,
    \top_I.branch[4].l_um_iw[103] ,
    \top_I.branch[4].l_um_iw[102] ,
    \top_I.branch[4].l_um_iw[101] ,
    \top_I.branch[4].l_um_iw[100] }),
    .uio_oe({\top_I.branch[4].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[4].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[4].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[0] }));
 tt_um_urish_dffram \top_I.branch[4].col_um[4].um_top_I.block_5_4.tt_um_I  (.clk(\top_I.branch[4].l_um_iw[162] ),
    .ena(\top_I.branch[4].l_um_ena[9] ),
    .rst_n(\top_I.branch[4].l_um_iw[163] ),
    .ui_in({\top_I.branch[4].l_um_iw[171] ,
    \top_I.branch[4].l_um_iw[170] ,
    \top_I.branch[4].l_um_iw[169] ,
    \top_I.branch[4].l_um_iw[168] ,
    \top_I.branch[4].l_um_iw[167] ,
    \top_I.branch[4].l_um_iw[166] ,
    \top_I.branch[4].l_um_iw[165] ,
    \top_I.branch[4].l_um_iw[164] }),
    .uio_in({\top_I.branch[4].l_um_iw[179] ,
    \top_I.branch[4].l_um_iw[178] ,
    \top_I.branch[4].l_um_iw[177] ,
    \top_I.branch[4].l_um_iw[176] ,
    \top_I.branch[4].l_um_iw[175] ,
    \top_I.branch[4].l_um_iw[174] ,
    \top_I.branch[4].l_um_iw[173] ,
    \top_I.branch[4].l_um_iw[172] }),
    .uio_oe({\top_I.branch[4].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[4].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[4].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[4].mux_I  (.k_one(\top_I.branch[4].l_k_one ),
    .k_zero(\top_I.branch[4].l_k_zero ),
    .addr({\top_I.branch[4].l_k_zero ,
    \top_I.branch[4].l_k_zero ,
    \top_I.branch[4].l_k_one ,
    \top_I.branch[4].l_k_zero ,
    \top_I.branch[4].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[4].l_um_ena[15] ,
    \top_I.branch[4].l_um_ena[14] ,
    \top_I.branch[4].l_um_ena[13] ,
    \top_I.branch[4].l_um_ena[12] ,
    \top_I.branch[4].l_um_ena[11] ,
    \top_I.branch[4].l_um_ena[10] ,
    \top_I.branch[4].l_um_ena[9] ,
    \top_I.branch[4].l_um_ena[8] ,
    \top_I.branch[4].l_um_ena[7] ,
    \top_I.branch[4].l_um_ena[6] ,
    \top_I.branch[4].l_um_ena[5] ,
    \top_I.branch[4].l_um_ena[4] ,
    \top_I.branch[4].l_um_ena[3] ,
    \top_I.branch[4].l_um_ena[2] ,
    \top_I.branch[4].l_um_ena[1] ,
    \top_I.branch[4].l_um_ena[0] }),
    .um_iw({\top_I.branch[4].l_um_iw[287] ,
    \top_I.branch[4].l_um_iw[286] ,
    \top_I.branch[4].l_um_iw[285] ,
    \top_I.branch[4].l_um_iw[284] ,
    \top_I.branch[4].l_um_iw[283] ,
    \top_I.branch[4].l_um_iw[282] ,
    \top_I.branch[4].l_um_iw[281] ,
    \top_I.branch[4].l_um_iw[280] ,
    \top_I.branch[4].l_um_iw[279] ,
    \top_I.branch[4].l_um_iw[278] ,
    \top_I.branch[4].l_um_iw[277] ,
    \top_I.branch[4].l_um_iw[276] ,
    \top_I.branch[4].l_um_iw[275] ,
    \top_I.branch[4].l_um_iw[274] ,
    \top_I.branch[4].l_um_iw[273] ,
    \top_I.branch[4].l_um_iw[272] ,
    \top_I.branch[4].l_um_iw[271] ,
    \top_I.branch[4].l_um_iw[270] ,
    \top_I.branch[4].l_um_iw[269] ,
    \top_I.branch[4].l_um_iw[268] ,
    \top_I.branch[4].l_um_iw[267] ,
    \top_I.branch[4].l_um_iw[266] ,
    \top_I.branch[4].l_um_iw[265] ,
    \top_I.branch[4].l_um_iw[264] ,
    \top_I.branch[4].l_um_iw[263] ,
    \top_I.branch[4].l_um_iw[262] ,
    \top_I.branch[4].l_um_iw[261] ,
    \top_I.branch[4].l_um_iw[260] ,
    \top_I.branch[4].l_um_iw[259] ,
    \top_I.branch[4].l_um_iw[258] ,
    \top_I.branch[4].l_um_iw[257] ,
    \top_I.branch[4].l_um_iw[256] ,
    \top_I.branch[4].l_um_iw[255] ,
    \top_I.branch[4].l_um_iw[254] ,
    \top_I.branch[4].l_um_iw[253] ,
    \top_I.branch[4].l_um_iw[252] ,
    \top_I.branch[4].l_um_iw[251] ,
    \top_I.branch[4].l_um_iw[250] ,
    \top_I.branch[4].l_um_iw[249] ,
    \top_I.branch[4].l_um_iw[248] ,
    \top_I.branch[4].l_um_iw[247] ,
    \top_I.branch[4].l_um_iw[246] ,
    \top_I.branch[4].l_um_iw[245] ,
    \top_I.branch[4].l_um_iw[244] ,
    \top_I.branch[4].l_um_iw[243] ,
    \top_I.branch[4].l_um_iw[242] ,
    \top_I.branch[4].l_um_iw[241] ,
    \top_I.branch[4].l_um_iw[240] ,
    \top_I.branch[4].l_um_iw[239] ,
    \top_I.branch[4].l_um_iw[238] ,
    \top_I.branch[4].l_um_iw[237] ,
    \top_I.branch[4].l_um_iw[236] ,
    \top_I.branch[4].l_um_iw[235] ,
    \top_I.branch[4].l_um_iw[234] ,
    \top_I.branch[4].l_um_iw[233] ,
    \top_I.branch[4].l_um_iw[232] ,
    \top_I.branch[4].l_um_iw[231] ,
    \top_I.branch[4].l_um_iw[230] ,
    \top_I.branch[4].l_um_iw[229] ,
    \top_I.branch[4].l_um_iw[228] ,
    \top_I.branch[4].l_um_iw[227] ,
    \top_I.branch[4].l_um_iw[226] ,
    \top_I.branch[4].l_um_iw[225] ,
    \top_I.branch[4].l_um_iw[224] ,
    \top_I.branch[4].l_um_iw[223] ,
    \top_I.branch[4].l_um_iw[222] ,
    \top_I.branch[4].l_um_iw[221] ,
    \top_I.branch[4].l_um_iw[220] ,
    \top_I.branch[4].l_um_iw[219] ,
    \top_I.branch[4].l_um_iw[218] ,
    \top_I.branch[4].l_um_iw[217] ,
    \top_I.branch[4].l_um_iw[216] ,
    \top_I.branch[4].l_um_iw[215] ,
    \top_I.branch[4].l_um_iw[214] ,
    \top_I.branch[4].l_um_iw[213] ,
    \top_I.branch[4].l_um_iw[212] ,
    \top_I.branch[4].l_um_iw[211] ,
    \top_I.branch[4].l_um_iw[210] ,
    \top_I.branch[4].l_um_iw[209] ,
    \top_I.branch[4].l_um_iw[208] ,
    \top_I.branch[4].l_um_iw[207] ,
    \top_I.branch[4].l_um_iw[206] ,
    \top_I.branch[4].l_um_iw[205] ,
    \top_I.branch[4].l_um_iw[204] ,
    \top_I.branch[4].l_um_iw[203] ,
    \top_I.branch[4].l_um_iw[202] ,
    \top_I.branch[4].l_um_iw[201] ,
    \top_I.branch[4].l_um_iw[200] ,
    \top_I.branch[4].l_um_iw[199] ,
    \top_I.branch[4].l_um_iw[198] ,
    \top_I.branch[4].l_um_iw[197] ,
    \top_I.branch[4].l_um_iw[196] ,
    \top_I.branch[4].l_um_iw[195] ,
    \top_I.branch[4].l_um_iw[194] ,
    \top_I.branch[4].l_um_iw[193] ,
    \top_I.branch[4].l_um_iw[192] ,
    \top_I.branch[4].l_um_iw[191] ,
    \top_I.branch[4].l_um_iw[190] ,
    \top_I.branch[4].l_um_iw[189] ,
    \top_I.branch[4].l_um_iw[188] ,
    \top_I.branch[4].l_um_iw[187] ,
    \top_I.branch[4].l_um_iw[186] ,
    \top_I.branch[4].l_um_iw[185] ,
    \top_I.branch[4].l_um_iw[184] ,
    \top_I.branch[4].l_um_iw[183] ,
    \top_I.branch[4].l_um_iw[182] ,
    \top_I.branch[4].l_um_iw[181] ,
    \top_I.branch[4].l_um_iw[180] ,
    \top_I.branch[4].l_um_iw[179] ,
    \top_I.branch[4].l_um_iw[178] ,
    \top_I.branch[4].l_um_iw[177] ,
    \top_I.branch[4].l_um_iw[176] ,
    \top_I.branch[4].l_um_iw[175] ,
    \top_I.branch[4].l_um_iw[174] ,
    \top_I.branch[4].l_um_iw[173] ,
    \top_I.branch[4].l_um_iw[172] ,
    \top_I.branch[4].l_um_iw[171] ,
    \top_I.branch[4].l_um_iw[170] ,
    \top_I.branch[4].l_um_iw[169] ,
    \top_I.branch[4].l_um_iw[168] ,
    \top_I.branch[4].l_um_iw[167] ,
    \top_I.branch[4].l_um_iw[166] ,
    \top_I.branch[4].l_um_iw[165] ,
    \top_I.branch[4].l_um_iw[164] ,
    \top_I.branch[4].l_um_iw[163] ,
    \top_I.branch[4].l_um_iw[162] ,
    \top_I.branch[4].l_um_iw[161] ,
    \top_I.branch[4].l_um_iw[160] ,
    \top_I.branch[4].l_um_iw[159] ,
    \top_I.branch[4].l_um_iw[158] ,
    \top_I.branch[4].l_um_iw[157] ,
    \top_I.branch[4].l_um_iw[156] ,
    \top_I.branch[4].l_um_iw[155] ,
    \top_I.branch[4].l_um_iw[154] ,
    \top_I.branch[4].l_um_iw[153] ,
    \top_I.branch[4].l_um_iw[152] ,
    \top_I.branch[4].l_um_iw[151] ,
    \top_I.branch[4].l_um_iw[150] ,
    \top_I.branch[4].l_um_iw[149] ,
    \top_I.branch[4].l_um_iw[148] ,
    \top_I.branch[4].l_um_iw[147] ,
    \top_I.branch[4].l_um_iw[146] ,
    \top_I.branch[4].l_um_iw[145] ,
    \top_I.branch[4].l_um_iw[144] ,
    \top_I.branch[4].l_um_iw[143] ,
    \top_I.branch[4].l_um_iw[142] ,
    \top_I.branch[4].l_um_iw[141] ,
    \top_I.branch[4].l_um_iw[140] ,
    \top_I.branch[4].l_um_iw[139] ,
    \top_I.branch[4].l_um_iw[138] ,
    \top_I.branch[4].l_um_iw[137] ,
    \top_I.branch[4].l_um_iw[136] ,
    \top_I.branch[4].l_um_iw[135] ,
    \top_I.branch[4].l_um_iw[134] ,
    \top_I.branch[4].l_um_iw[133] ,
    \top_I.branch[4].l_um_iw[132] ,
    \top_I.branch[4].l_um_iw[131] ,
    \top_I.branch[4].l_um_iw[130] ,
    \top_I.branch[4].l_um_iw[129] ,
    \top_I.branch[4].l_um_iw[128] ,
    \top_I.branch[4].l_um_iw[127] ,
    \top_I.branch[4].l_um_iw[126] ,
    \top_I.branch[4].l_um_iw[125] ,
    \top_I.branch[4].l_um_iw[124] ,
    \top_I.branch[4].l_um_iw[123] ,
    \top_I.branch[4].l_um_iw[122] ,
    \top_I.branch[4].l_um_iw[121] ,
    \top_I.branch[4].l_um_iw[120] ,
    \top_I.branch[4].l_um_iw[119] ,
    \top_I.branch[4].l_um_iw[118] ,
    \top_I.branch[4].l_um_iw[117] ,
    \top_I.branch[4].l_um_iw[116] ,
    \top_I.branch[4].l_um_iw[115] ,
    \top_I.branch[4].l_um_iw[114] ,
    \top_I.branch[4].l_um_iw[113] ,
    \top_I.branch[4].l_um_iw[112] ,
    \top_I.branch[4].l_um_iw[111] ,
    \top_I.branch[4].l_um_iw[110] ,
    \top_I.branch[4].l_um_iw[109] ,
    \top_I.branch[4].l_um_iw[108] ,
    \top_I.branch[4].l_um_iw[107] ,
    \top_I.branch[4].l_um_iw[106] ,
    \top_I.branch[4].l_um_iw[105] ,
    \top_I.branch[4].l_um_iw[104] ,
    \top_I.branch[4].l_um_iw[103] ,
    \top_I.branch[4].l_um_iw[102] ,
    \top_I.branch[4].l_um_iw[101] ,
    \top_I.branch[4].l_um_iw[100] ,
    \top_I.branch[4].l_um_iw[99] ,
    \top_I.branch[4].l_um_iw[98] ,
    \top_I.branch[4].l_um_iw[97] ,
    \top_I.branch[4].l_um_iw[96] ,
    \top_I.branch[4].l_um_iw[95] ,
    \top_I.branch[4].l_um_iw[94] ,
    \top_I.branch[4].l_um_iw[93] ,
    \top_I.branch[4].l_um_iw[92] ,
    \top_I.branch[4].l_um_iw[91] ,
    \top_I.branch[4].l_um_iw[90] ,
    \top_I.branch[4].l_um_iw[89] ,
    \top_I.branch[4].l_um_iw[88] ,
    \top_I.branch[4].l_um_iw[87] ,
    \top_I.branch[4].l_um_iw[86] ,
    \top_I.branch[4].l_um_iw[85] ,
    \top_I.branch[4].l_um_iw[84] ,
    \top_I.branch[4].l_um_iw[83] ,
    \top_I.branch[4].l_um_iw[82] ,
    \top_I.branch[4].l_um_iw[81] ,
    \top_I.branch[4].l_um_iw[80] ,
    \top_I.branch[4].l_um_iw[79] ,
    \top_I.branch[4].l_um_iw[78] ,
    \top_I.branch[4].l_um_iw[77] ,
    \top_I.branch[4].l_um_iw[76] ,
    \top_I.branch[4].l_um_iw[75] ,
    \top_I.branch[4].l_um_iw[74] ,
    \top_I.branch[4].l_um_iw[73] ,
    \top_I.branch[4].l_um_iw[72] ,
    \top_I.branch[4].l_um_iw[71] ,
    \top_I.branch[4].l_um_iw[70] ,
    \top_I.branch[4].l_um_iw[69] ,
    \top_I.branch[4].l_um_iw[68] ,
    \top_I.branch[4].l_um_iw[67] ,
    \top_I.branch[4].l_um_iw[66] ,
    \top_I.branch[4].l_um_iw[65] ,
    \top_I.branch[4].l_um_iw[64] ,
    \top_I.branch[4].l_um_iw[63] ,
    \top_I.branch[4].l_um_iw[62] ,
    \top_I.branch[4].l_um_iw[61] ,
    \top_I.branch[4].l_um_iw[60] ,
    \top_I.branch[4].l_um_iw[59] ,
    \top_I.branch[4].l_um_iw[58] ,
    \top_I.branch[4].l_um_iw[57] ,
    \top_I.branch[4].l_um_iw[56] ,
    \top_I.branch[4].l_um_iw[55] ,
    \top_I.branch[4].l_um_iw[54] ,
    \top_I.branch[4].l_um_iw[53] ,
    \top_I.branch[4].l_um_iw[52] ,
    \top_I.branch[4].l_um_iw[51] ,
    \top_I.branch[4].l_um_iw[50] ,
    \top_I.branch[4].l_um_iw[49] ,
    \top_I.branch[4].l_um_iw[48] ,
    \top_I.branch[4].l_um_iw[47] ,
    \top_I.branch[4].l_um_iw[46] ,
    \top_I.branch[4].l_um_iw[45] ,
    \top_I.branch[4].l_um_iw[44] ,
    \top_I.branch[4].l_um_iw[43] ,
    \top_I.branch[4].l_um_iw[42] ,
    \top_I.branch[4].l_um_iw[41] ,
    \top_I.branch[4].l_um_iw[40] ,
    \top_I.branch[4].l_um_iw[39] ,
    \top_I.branch[4].l_um_iw[38] ,
    \top_I.branch[4].l_um_iw[37] ,
    \top_I.branch[4].l_um_iw[36] ,
    \top_I.branch[4].l_um_iw[35] ,
    \top_I.branch[4].l_um_iw[34] ,
    \top_I.branch[4].l_um_iw[33] ,
    \top_I.branch[4].l_um_iw[32] ,
    \top_I.branch[4].l_um_iw[31] ,
    \top_I.branch[4].l_um_iw[30] ,
    \top_I.branch[4].l_um_iw[29] ,
    \top_I.branch[4].l_um_iw[28] ,
    \top_I.branch[4].l_um_iw[27] ,
    \top_I.branch[4].l_um_iw[26] ,
    \top_I.branch[4].l_um_iw[25] ,
    \top_I.branch[4].l_um_iw[24] ,
    \top_I.branch[4].l_um_iw[23] ,
    \top_I.branch[4].l_um_iw[22] ,
    \top_I.branch[4].l_um_iw[21] ,
    \top_I.branch[4].l_um_iw[20] ,
    \top_I.branch[4].l_um_iw[19] ,
    \top_I.branch[4].l_um_iw[18] ,
    \top_I.branch[4].l_um_iw[17] ,
    \top_I.branch[4].l_um_iw[16] ,
    \top_I.branch[4].l_um_iw[15] ,
    \top_I.branch[4].l_um_iw[14] ,
    \top_I.branch[4].l_um_iw[13] ,
    \top_I.branch[4].l_um_iw[12] ,
    \top_I.branch[4].l_um_iw[11] ,
    \top_I.branch[4].l_um_iw[10] ,
    \top_I.branch[4].l_um_iw[9] ,
    \top_I.branch[4].l_um_iw[8] ,
    \top_I.branch[4].l_um_iw[7] ,
    \top_I.branch[4].l_um_iw[6] ,
    \top_I.branch[4].l_um_iw[5] ,
    \top_I.branch[4].l_um_iw[4] ,
    \top_I.branch[4].l_um_iw[3] ,
    \top_I.branch[4].l_um_iw[2] ,
    \top_I.branch[4].l_um_iw[1] ,
    \top_I.branch[4].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[9] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[5] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[15] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[14] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[13] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[12] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[11] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].l_um_k_zero[10] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_oe[0] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uio_out[0] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[7] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[6] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[5] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[4] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[3] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[2] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[1] ,
    \top_I.branch[4].col_um[4].um_top_I.uo_out[0] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[8] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[7] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].l_um_k_zero[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_oe[0] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uio_out[0] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[7] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[6] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[5] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[4] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[3] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[2] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[1] ,
    \top_I.branch[4].col_um[2].um_top_I.uo_out[0] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[4] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[3] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[2] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].l_um_k_zero[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[4].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[5].col_um[0].um_bot_I.block_4_16.tt_um_I  (.clk(\top_I.branch[5].l_um_iw[0] ),
    .ena(\top_I.branch[5].l_um_ena[0] ),
    .rst_n(\top_I.branch[5].l_um_iw[1] ),
    .ui_in({\top_I.branch[5].l_um_iw[9] ,
    \top_I.branch[5].l_um_iw[8] ,
    \top_I.branch[5].l_um_iw[7] ,
    \top_I.branch[5].l_um_iw[6] ,
    \top_I.branch[5].l_um_iw[5] ,
    \top_I.branch[5].l_um_iw[4] ,
    \top_I.branch[5].l_um_iw[3] ,
    \top_I.branch[5].l_um_iw[2] }),
    .uio_in({\top_I.branch[5].l_um_iw[17] ,
    \top_I.branch[5].l_um_iw[16] ,
    \top_I.branch[5].l_um_iw[15] ,
    \top_I.branch[5].l_um_iw[14] ,
    \top_I.branch[5].l_um_iw[13] ,
    \top_I.branch[5].l_um_iw[12] ,
    \top_I.branch[5].l_um_iw[11] ,
    \top_I.branch[5].l_um_iw[10] }),
    .uio_oe({\top_I.branch[5].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[5].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[5].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[5].mux_I  (.k_one(\top_I.branch[5].l_k_one ),
    .k_zero(\top_I.branch[5].l_k_zero ),
    .addr({\top_I.branch[5].l_k_zero ,
    \top_I.branch[5].l_k_zero ,
    \top_I.branch[5].l_k_one ,
    \top_I.branch[5].l_k_zero ,
    \top_I.branch[5].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[5].l_um_ena[15] ,
    \top_I.branch[5].l_um_ena[14] ,
    \top_I.branch[5].l_um_ena[13] ,
    \top_I.branch[5].l_um_ena[12] ,
    \top_I.branch[5].l_um_ena[11] ,
    \top_I.branch[5].l_um_ena[10] ,
    \top_I.branch[5].l_um_ena[9] ,
    \top_I.branch[5].l_um_ena[8] ,
    \top_I.branch[5].l_um_ena[7] ,
    \top_I.branch[5].l_um_ena[6] ,
    \top_I.branch[5].l_um_ena[5] ,
    \top_I.branch[5].l_um_ena[4] ,
    \top_I.branch[5].l_um_ena[3] ,
    \top_I.branch[5].l_um_ena[2] ,
    \top_I.branch[5].l_um_ena[1] ,
    \top_I.branch[5].l_um_ena[0] }),
    .um_iw({\top_I.branch[5].l_um_iw[287] ,
    \top_I.branch[5].l_um_iw[286] ,
    \top_I.branch[5].l_um_iw[285] ,
    \top_I.branch[5].l_um_iw[284] ,
    \top_I.branch[5].l_um_iw[283] ,
    \top_I.branch[5].l_um_iw[282] ,
    \top_I.branch[5].l_um_iw[281] ,
    \top_I.branch[5].l_um_iw[280] ,
    \top_I.branch[5].l_um_iw[279] ,
    \top_I.branch[5].l_um_iw[278] ,
    \top_I.branch[5].l_um_iw[277] ,
    \top_I.branch[5].l_um_iw[276] ,
    \top_I.branch[5].l_um_iw[275] ,
    \top_I.branch[5].l_um_iw[274] ,
    \top_I.branch[5].l_um_iw[273] ,
    \top_I.branch[5].l_um_iw[272] ,
    \top_I.branch[5].l_um_iw[271] ,
    \top_I.branch[5].l_um_iw[270] ,
    \top_I.branch[5].l_um_iw[269] ,
    \top_I.branch[5].l_um_iw[268] ,
    \top_I.branch[5].l_um_iw[267] ,
    \top_I.branch[5].l_um_iw[266] ,
    \top_I.branch[5].l_um_iw[265] ,
    \top_I.branch[5].l_um_iw[264] ,
    \top_I.branch[5].l_um_iw[263] ,
    \top_I.branch[5].l_um_iw[262] ,
    \top_I.branch[5].l_um_iw[261] ,
    \top_I.branch[5].l_um_iw[260] ,
    \top_I.branch[5].l_um_iw[259] ,
    \top_I.branch[5].l_um_iw[258] ,
    \top_I.branch[5].l_um_iw[257] ,
    \top_I.branch[5].l_um_iw[256] ,
    \top_I.branch[5].l_um_iw[255] ,
    \top_I.branch[5].l_um_iw[254] ,
    \top_I.branch[5].l_um_iw[253] ,
    \top_I.branch[5].l_um_iw[252] ,
    \top_I.branch[5].l_um_iw[251] ,
    \top_I.branch[5].l_um_iw[250] ,
    \top_I.branch[5].l_um_iw[249] ,
    \top_I.branch[5].l_um_iw[248] ,
    \top_I.branch[5].l_um_iw[247] ,
    \top_I.branch[5].l_um_iw[246] ,
    \top_I.branch[5].l_um_iw[245] ,
    \top_I.branch[5].l_um_iw[244] ,
    \top_I.branch[5].l_um_iw[243] ,
    \top_I.branch[5].l_um_iw[242] ,
    \top_I.branch[5].l_um_iw[241] ,
    \top_I.branch[5].l_um_iw[240] ,
    \top_I.branch[5].l_um_iw[239] ,
    \top_I.branch[5].l_um_iw[238] ,
    \top_I.branch[5].l_um_iw[237] ,
    \top_I.branch[5].l_um_iw[236] ,
    \top_I.branch[5].l_um_iw[235] ,
    \top_I.branch[5].l_um_iw[234] ,
    \top_I.branch[5].l_um_iw[233] ,
    \top_I.branch[5].l_um_iw[232] ,
    \top_I.branch[5].l_um_iw[231] ,
    \top_I.branch[5].l_um_iw[230] ,
    \top_I.branch[5].l_um_iw[229] ,
    \top_I.branch[5].l_um_iw[228] ,
    \top_I.branch[5].l_um_iw[227] ,
    \top_I.branch[5].l_um_iw[226] ,
    \top_I.branch[5].l_um_iw[225] ,
    \top_I.branch[5].l_um_iw[224] ,
    \top_I.branch[5].l_um_iw[223] ,
    \top_I.branch[5].l_um_iw[222] ,
    \top_I.branch[5].l_um_iw[221] ,
    \top_I.branch[5].l_um_iw[220] ,
    \top_I.branch[5].l_um_iw[219] ,
    \top_I.branch[5].l_um_iw[218] ,
    \top_I.branch[5].l_um_iw[217] ,
    \top_I.branch[5].l_um_iw[216] ,
    \top_I.branch[5].l_um_iw[215] ,
    \top_I.branch[5].l_um_iw[214] ,
    \top_I.branch[5].l_um_iw[213] ,
    \top_I.branch[5].l_um_iw[212] ,
    \top_I.branch[5].l_um_iw[211] ,
    \top_I.branch[5].l_um_iw[210] ,
    \top_I.branch[5].l_um_iw[209] ,
    \top_I.branch[5].l_um_iw[208] ,
    \top_I.branch[5].l_um_iw[207] ,
    \top_I.branch[5].l_um_iw[206] ,
    \top_I.branch[5].l_um_iw[205] ,
    \top_I.branch[5].l_um_iw[204] ,
    \top_I.branch[5].l_um_iw[203] ,
    \top_I.branch[5].l_um_iw[202] ,
    \top_I.branch[5].l_um_iw[201] ,
    \top_I.branch[5].l_um_iw[200] ,
    \top_I.branch[5].l_um_iw[199] ,
    \top_I.branch[5].l_um_iw[198] ,
    \top_I.branch[5].l_um_iw[197] ,
    \top_I.branch[5].l_um_iw[196] ,
    \top_I.branch[5].l_um_iw[195] ,
    \top_I.branch[5].l_um_iw[194] ,
    \top_I.branch[5].l_um_iw[193] ,
    \top_I.branch[5].l_um_iw[192] ,
    \top_I.branch[5].l_um_iw[191] ,
    \top_I.branch[5].l_um_iw[190] ,
    \top_I.branch[5].l_um_iw[189] ,
    \top_I.branch[5].l_um_iw[188] ,
    \top_I.branch[5].l_um_iw[187] ,
    \top_I.branch[5].l_um_iw[186] ,
    \top_I.branch[5].l_um_iw[185] ,
    \top_I.branch[5].l_um_iw[184] ,
    \top_I.branch[5].l_um_iw[183] ,
    \top_I.branch[5].l_um_iw[182] ,
    \top_I.branch[5].l_um_iw[181] ,
    \top_I.branch[5].l_um_iw[180] ,
    \top_I.branch[5].l_um_iw[179] ,
    \top_I.branch[5].l_um_iw[178] ,
    \top_I.branch[5].l_um_iw[177] ,
    \top_I.branch[5].l_um_iw[176] ,
    \top_I.branch[5].l_um_iw[175] ,
    \top_I.branch[5].l_um_iw[174] ,
    \top_I.branch[5].l_um_iw[173] ,
    \top_I.branch[5].l_um_iw[172] ,
    \top_I.branch[5].l_um_iw[171] ,
    \top_I.branch[5].l_um_iw[170] ,
    \top_I.branch[5].l_um_iw[169] ,
    \top_I.branch[5].l_um_iw[168] ,
    \top_I.branch[5].l_um_iw[167] ,
    \top_I.branch[5].l_um_iw[166] ,
    \top_I.branch[5].l_um_iw[165] ,
    \top_I.branch[5].l_um_iw[164] ,
    \top_I.branch[5].l_um_iw[163] ,
    \top_I.branch[5].l_um_iw[162] ,
    \top_I.branch[5].l_um_iw[161] ,
    \top_I.branch[5].l_um_iw[160] ,
    \top_I.branch[5].l_um_iw[159] ,
    \top_I.branch[5].l_um_iw[158] ,
    \top_I.branch[5].l_um_iw[157] ,
    \top_I.branch[5].l_um_iw[156] ,
    \top_I.branch[5].l_um_iw[155] ,
    \top_I.branch[5].l_um_iw[154] ,
    \top_I.branch[5].l_um_iw[153] ,
    \top_I.branch[5].l_um_iw[152] ,
    \top_I.branch[5].l_um_iw[151] ,
    \top_I.branch[5].l_um_iw[150] ,
    \top_I.branch[5].l_um_iw[149] ,
    \top_I.branch[5].l_um_iw[148] ,
    \top_I.branch[5].l_um_iw[147] ,
    \top_I.branch[5].l_um_iw[146] ,
    \top_I.branch[5].l_um_iw[145] ,
    \top_I.branch[5].l_um_iw[144] ,
    \top_I.branch[5].l_um_iw[143] ,
    \top_I.branch[5].l_um_iw[142] ,
    \top_I.branch[5].l_um_iw[141] ,
    \top_I.branch[5].l_um_iw[140] ,
    \top_I.branch[5].l_um_iw[139] ,
    \top_I.branch[5].l_um_iw[138] ,
    \top_I.branch[5].l_um_iw[137] ,
    \top_I.branch[5].l_um_iw[136] ,
    \top_I.branch[5].l_um_iw[135] ,
    \top_I.branch[5].l_um_iw[134] ,
    \top_I.branch[5].l_um_iw[133] ,
    \top_I.branch[5].l_um_iw[132] ,
    \top_I.branch[5].l_um_iw[131] ,
    \top_I.branch[5].l_um_iw[130] ,
    \top_I.branch[5].l_um_iw[129] ,
    \top_I.branch[5].l_um_iw[128] ,
    \top_I.branch[5].l_um_iw[127] ,
    \top_I.branch[5].l_um_iw[126] ,
    \top_I.branch[5].l_um_iw[125] ,
    \top_I.branch[5].l_um_iw[124] ,
    \top_I.branch[5].l_um_iw[123] ,
    \top_I.branch[5].l_um_iw[122] ,
    \top_I.branch[5].l_um_iw[121] ,
    \top_I.branch[5].l_um_iw[120] ,
    \top_I.branch[5].l_um_iw[119] ,
    \top_I.branch[5].l_um_iw[118] ,
    \top_I.branch[5].l_um_iw[117] ,
    \top_I.branch[5].l_um_iw[116] ,
    \top_I.branch[5].l_um_iw[115] ,
    \top_I.branch[5].l_um_iw[114] ,
    \top_I.branch[5].l_um_iw[113] ,
    \top_I.branch[5].l_um_iw[112] ,
    \top_I.branch[5].l_um_iw[111] ,
    \top_I.branch[5].l_um_iw[110] ,
    \top_I.branch[5].l_um_iw[109] ,
    \top_I.branch[5].l_um_iw[108] ,
    \top_I.branch[5].l_um_iw[107] ,
    \top_I.branch[5].l_um_iw[106] ,
    \top_I.branch[5].l_um_iw[105] ,
    \top_I.branch[5].l_um_iw[104] ,
    \top_I.branch[5].l_um_iw[103] ,
    \top_I.branch[5].l_um_iw[102] ,
    \top_I.branch[5].l_um_iw[101] ,
    \top_I.branch[5].l_um_iw[100] ,
    \top_I.branch[5].l_um_iw[99] ,
    \top_I.branch[5].l_um_iw[98] ,
    \top_I.branch[5].l_um_iw[97] ,
    \top_I.branch[5].l_um_iw[96] ,
    \top_I.branch[5].l_um_iw[95] ,
    \top_I.branch[5].l_um_iw[94] ,
    \top_I.branch[5].l_um_iw[93] ,
    \top_I.branch[5].l_um_iw[92] ,
    \top_I.branch[5].l_um_iw[91] ,
    \top_I.branch[5].l_um_iw[90] ,
    \top_I.branch[5].l_um_iw[89] ,
    \top_I.branch[5].l_um_iw[88] ,
    \top_I.branch[5].l_um_iw[87] ,
    \top_I.branch[5].l_um_iw[86] ,
    \top_I.branch[5].l_um_iw[85] ,
    \top_I.branch[5].l_um_iw[84] ,
    \top_I.branch[5].l_um_iw[83] ,
    \top_I.branch[5].l_um_iw[82] ,
    \top_I.branch[5].l_um_iw[81] ,
    \top_I.branch[5].l_um_iw[80] ,
    \top_I.branch[5].l_um_iw[79] ,
    \top_I.branch[5].l_um_iw[78] ,
    \top_I.branch[5].l_um_iw[77] ,
    \top_I.branch[5].l_um_iw[76] ,
    \top_I.branch[5].l_um_iw[75] ,
    \top_I.branch[5].l_um_iw[74] ,
    \top_I.branch[5].l_um_iw[73] ,
    \top_I.branch[5].l_um_iw[72] ,
    \top_I.branch[5].l_um_iw[71] ,
    \top_I.branch[5].l_um_iw[70] ,
    \top_I.branch[5].l_um_iw[69] ,
    \top_I.branch[5].l_um_iw[68] ,
    \top_I.branch[5].l_um_iw[67] ,
    \top_I.branch[5].l_um_iw[66] ,
    \top_I.branch[5].l_um_iw[65] ,
    \top_I.branch[5].l_um_iw[64] ,
    \top_I.branch[5].l_um_iw[63] ,
    \top_I.branch[5].l_um_iw[62] ,
    \top_I.branch[5].l_um_iw[61] ,
    \top_I.branch[5].l_um_iw[60] ,
    \top_I.branch[5].l_um_iw[59] ,
    \top_I.branch[5].l_um_iw[58] ,
    \top_I.branch[5].l_um_iw[57] ,
    \top_I.branch[5].l_um_iw[56] ,
    \top_I.branch[5].l_um_iw[55] ,
    \top_I.branch[5].l_um_iw[54] ,
    \top_I.branch[5].l_um_iw[53] ,
    \top_I.branch[5].l_um_iw[52] ,
    \top_I.branch[5].l_um_iw[51] ,
    \top_I.branch[5].l_um_iw[50] ,
    \top_I.branch[5].l_um_iw[49] ,
    \top_I.branch[5].l_um_iw[48] ,
    \top_I.branch[5].l_um_iw[47] ,
    \top_I.branch[5].l_um_iw[46] ,
    \top_I.branch[5].l_um_iw[45] ,
    \top_I.branch[5].l_um_iw[44] ,
    \top_I.branch[5].l_um_iw[43] ,
    \top_I.branch[5].l_um_iw[42] ,
    \top_I.branch[5].l_um_iw[41] ,
    \top_I.branch[5].l_um_iw[40] ,
    \top_I.branch[5].l_um_iw[39] ,
    \top_I.branch[5].l_um_iw[38] ,
    \top_I.branch[5].l_um_iw[37] ,
    \top_I.branch[5].l_um_iw[36] ,
    \top_I.branch[5].l_um_iw[35] ,
    \top_I.branch[5].l_um_iw[34] ,
    \top_I.branch[5].l_um_iw[33] ,
    \top_I.branch[5].l_um_iw[32] ,
    \top_I.branch[5].l_um_iw[31] ,
    \top_I.branch[5].l_um_iw[30] ,
    \top_I.branch[5].l_um_iw[29] ,
    \top_I.branch[5].l_um_iw[28] ,
    \top_I.branch[5].l_um_iw[27] ,
    \top_I.branch[5].l_um_iw[26] ,
    \top_I.branch[5].l_um_iw[25] ,
    \top_I.branch[5].l_um_iw[24] ,
    \top_I.branch[5].l_um_iw[23] ,
    \top_I.branch[5].l_um_iw[22] ,
    \top_I.branch[5].l_um_iw[21] ,
    \top_I.branch[5].l_um_iw[20] ,
    \top_I.branch[5].l_um_iw[19] ,
    \top_I.branch[5].l_um_iw[18] ,
    \top_I.branch[5].l_um_iw[17] ,
    \top_I.branch[5].l_um_iw[16] ,
    \top_I.branch[5].l_um_iw[15] ,
    \top_I.branch[5].l_um_iw[14] ,
    \top_I.branch[5].l_um_iw[13] ,
    \top_I.branch[5].l_um_iw[12] ,
    \top_I.branch[5].l_um_iw[11] ,
    \top_I.branch[5].l_um_iw[10] ,
    \top_I.branch[5].l_um_iw[9] ,
    \top_I.branch[5].l_um_iw[8] ,
    \top_I.branch[5].l_um_iw[7] ,
    \top_I.branch[5].l_um_iw[6] ,
    \top_I.branch[5].l_um_iw[5] ,
    \top_I.branch[5].l_um_iw[4] ,
    \top_I.branch[5].l_um_iw[3] ,
    \top_I.branch[5].l_um_iw[2] ,
    \top_I.branch[5].l_um_iw[1] ,
    \top_I.branch[5].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[15] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[14] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[13] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[12] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[11] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[10] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[9] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[8] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[7] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[6] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[5] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[4] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[3] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[2] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].l_um_k_zero[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[5].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[6].col_um[0].um_top_I.block_7_0.tt_um_I  (.clk(\top_I.branch[6].l_um_iw[18] ),
    .ena(\top_I.branch[6].l_um_ena[1] ),
    .rst_n(\top_I.branch[6].l_um_iw[19] ),
    .ui_in({\top_I.branch[6].l_um_iw[27] ,
    \top_I.branch[6].l_um_iw[26] ,
    \top_I.branch[6].l_um_iw[25] ,
    \top_I.branch[6].l_um_iw[24] ,
    \top_I.branch[6].l_um_iw[23] ,
    \top_I.branch[6].l_um_iw[22] ,
    \top_I.branch[6].l_um_iw[21] ,
    \top_I.branch[6].l_um_iw[20] }),
    .uio_in({\top_I.branch[6].l_um_iw[35] ,
    \top_I.branch[6].l_um_iw[34] ,
    \top_I.branch[6].l_um_iw[33] ,
    \top_I.branch[6].l_um_iw[32] ,
    \top_I.branch[6].l_um_iw[31] ,
    \top_I.branch[6].l_um_iw[30] ,
    \top_I.branch[6].l_um_iw[29] ,
    \top_I.branch[6].l_um_iw[28] }),
    .uio_oe({\top_I.branch[6].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[6].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[6].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[6].mux_I  (.k_one(\top_I.branch[6].l_k_one ),
    .k_zero(\top_I.branch[6].l_k_zero ),
    .addr({\top_I.branch[6].l_k_zero ,
    \top_I.branch[6].l_k_zero ,
    \top_I.branch[6].l_k_one ,
    \top_I.branch[6].l_k_one ,
    \top_I.branch[6].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[6].l_um_ena[15] ,
    \top_I.branch[6].l_um_ena[14] ,
    \top_I.branch[6].l_um_ena[13] ,
    \top_I.branch[6].l_um_ena[12] ,
    \top_I.branch[6].l_um_ena[11] ,
    \top_I.branch[6].l_um_ena[10] ,
    \top_I.branch[6].l_um_ena[9] ,
    \top_I.branch[6].l_um_ena[8] ,
    \top_I.branch[6].l_um_ena[7] ,
    \top_I.branch[6].l_um_ena[6] ,
    \top_I.branch[6].l_um_ena[5] ,
    \top_I.branch[6].l_um_ena[4] ,
    \top_I.branch[6].l_um_ena[3] ,
    \top_I.branch[6].l_um_ena[2] ,
    \top_I.branch[6].l_um_ena[1] ,
    \top_I.branch[6].l_um_ena[0] }),
    .um_iw({\top_I.branch[6].l_um_iw[287] ,
    \top_I.branch[6].l_um_iw[286] ,
    \top_I.branch[6].l_um_iw[285] ,
    \top_I.branch[6].l_um_iw[284] ,
    \top_I.branch[6].l_um_iw[283] ,
    \top_I.branch[6].l_um_iw[282] ,
    \top_I.branch[6].l_um_iw[281] ,
    \top_I.branch[6].l_um_iw[280] ,
    \top_I.branch[6].l_um_iw[279] ,
    \top_I.branch[6].l_um_iw[278] ,
    \top_I.branch[6].l_um_iw[277] ,
    \top_I.branch[6].l_um_iw[276] ,
    \top_I.branch[6].l_um_iw[275] ,
    \top_I.branch[6].l_um_iw[274] ,
    \top_I.branch[6].l_um_iw[273] ,
    \top_I.branch[6].l_um_iw[272] ,
    \top_I.branch[6].l_um_iw[271] ,
    \top_I.branch[6].l_um_iw[270] ,
    \top_I.branch[6].l_um_iw[269] ,
    \top_I.branch[6].l_um_iw[268] ,
    \top_I.branch[6].l_um_iw[267] ,
    \top_I.branch[6].l_um_iw[266] ,
    \top_I.branch[6].l_um_iw[265] ,
    \top_I.branch[6].l_um_iw[264] ,
    \top_I.branch[6].l_um_iw[263] ,
    \top_I.branch[6].l_um_iw[262] ,
    \top_I.branch[6].l_um_iw[261] ,
    \top_I.branch[6].l_um_iw[260] ,
    \top_I.branch[6].l_um_iw[259] ,
    \top_I.branch[6].l_um_iw[258] ,
    \top_I.branch[6].l_um_iw[257] ,
    \top_I.branch[6].l_um_iw[256] ,
    \top_I.branch[6].l_um_iw[255] ,
    \top_I.branch[6].l_um_iw[254] ,
    \top_I.branch[6].l_um_iw[253] ,
    \top_I.branch[6].l_um_iw[252] ,
    \top_I.branch[6].l_um_iw[251] ,
    \top_I.branch[6].l_um_iw[250] ,
    \top_I.branch[6].l_um_iw[249] ,
    \top_I.branch[6].l_um_iw[248] ,
    \top_I.branch[6].l_um_iw[247] ,
    \top_I.branch[6].l_um_iw[246] ,
    \top_I.branch[6].l_um_iw[245] ,
    \top_I.branch[6].l_um_iw[244] ,
    \top_I.branch[6].l_um_iw[243] ,
    \top_I.branch[6].l_um_iw[242] ,
    \top_I.branch[6].l_um_iw[241] ,
    \top_I.branch[6].l_um_iw[240] ,
    \top_I.branch[6].l_um_iw[239] ,
    \top_I.branch[6].l_um_iw[238] ,
    \top_I.branch[6].l_um_iw[237] ,
    \top_I.branch[6].l_um_iw[236] ,
    \top_I.branch[6].l_um_iw[235] ,
    \top_I.branch[6].l_um_iw[234] ,
    \top_I.branch[6].l_um_iw[233] ,
    \top_I.branch[6].l_um_iw[232] ,
    \top_I.branch[6].l_um_iw[231] ,
    \top_I.branch[6].l_um_iw[230] ,
    \top_I.branch[6].l_um_iw[229] ,
    \top_I.branch[6].l_um_iw[228] ,
    \top_I.branch[6].l_um_iw[227] ,
    \top_I.branch[6].l_um_iw[226] ,
    \top_I.branch[6].l_um_iw[225] ,
    \top_I.branch[6].l_um_iw[224] ,
    \top_I.branch[6].l_um_iw[223] ,
    \top_I.branch[6].l_um_iw[222] ,
    \top_I.branch[6].l_um_iw[221] ,
    \top_I.branch[6].l_um_iw[220] ,
    \top_I.branch[6].l_um_iw[219] ,
    \top_I.branch[6].l_um_iw[218] ,
    \top_I.branch[6].l_um_iw[217] ,
    \top_I.branch[6].l_um_iw[216] ,
    \top_I.branch[6].l_um_iw[215] ,
    \top_I.branch[6].l_um_iw[214] ,
    \top_I.branch[6].l_um_iw[213] ,
    \top_I.branch[6].l_um_iw[212] ,
    \top_I.branch[6].l_um_iw[211] ,
    \top_I.branch[6].l_um_iw[210] ,
    \top_I.branch[6].l_um_iw[209] ,
    \top_I.branch[6].l_um_iw[208] ,
    \top_I.branch[6].l_um_iw[207] ,
    \top_I.branch[6].l_um_iw[206] ,
    \top_I.branch[6].l_um_iw[205] ,
    \top_I.branch[6].l_um_iw[204] ,
    \top_I.branch[6].l_um_iw[203] ,
    \top_I.branch[6].l_um_iw[202] ,
    \top_I.branch[6].l_um_iw[201] ,
    \top_I.branch[6].l_um_iw[200] ,
    \top_I.branch[6].l_um_iw[199] ,
    \top_I.branch[6].l_um_iw[198] ,
    \top_I.branch[6].l_um_iw[197] ,
    \top_I.branch[6].l_um_iw[196] ,
    \top_I.branch[6].l_um_iw[195] ,
    \top_I.branch[6].l_um_iw[194] ,
    \top_I.branch[6].l_um_iw[193] ,
    \top_I.branch[6].l_um_iw[192] ,
    \top_I.branch[6].l_um_iw[191] ,
    \top_I.branch[6].l_um_iw[190] ,
    \top_I.branch[6].l_um_iw[189] ,
    \top_I.branch[6].l_um_iw[188] ,
    \top_I.branch[6].l_um_iw[187] ,
    \top_I.branch[6].l_um_iw[186] ,
    \top_I.branch[6].l_um_iw[185] ,
    \top_I.branch[6].l_um_iw[184] ,
    \top_I.branch[6].l_um_iw[183] ,
    \top_I.branch[6].l_um_iw[182] ,
    \top_I.branch[6].l_um_iw[181] ,
    \top_I.branch[6].l_um_iw[180] ,
    \top_I.branch[6].l_um_iw[179] ,
    \top_I.branch[6].l_um_iw[178] ,
    \top_I.branch[6].l_um_iw[177] ,
    \top_I.branch[6].l_um_iw[176] ,
    \top_I.branch[6].l_um_iw[175] ,
    \top_I.branch[6].l_um_iw[174] ,
    \top_I.branch[6].l_um_iw[173] ,
    \top_I.branch[6].l_um_iw[172] ,
    \top_I.branch[6].l_um_iw[171] ,
    \top_I.branch[6].l_um_iw[170] ,
    \top_I.branch[6].l_um_iw[169] ,
    \top_I.branch[6].l_um_iw[168] ,
    \top_I.branch[6].l_um_iw[167] ,
    \top_I.branch[6].l_um_iw[166] ,
    \top_I.branch[6].l_um_iw[165] ,
    \top_I.branch[6].l_um_iw[164] ,
    \top_I.branch[6].l_um_iw[163] ,
    \top_I.branch[6].l_um_iw[162] ,
    \top_I.branch[6].l_um_iw[161] ,
    \top_I.branch[6].l_um_iw[160] ,
    \top_I.branch[6].l_um_iw[159] ,
    \top_I.branch[6].l_um_iw[158] ,
    \top_I.branch[6].l_um_iw[157] ,
    \top_I.branch[6].l_um_iw[156] ,
    \top_I.branch[6].l_um_iw[155] ,
    \top_I.branch[6].l_um_iw[154] ,
    \top_I.branch[6].l_um_iw[153] ,
    \top_I.branch[6].l_um_iw[152] ,
    \top_I.branch[6].l_um_iw[151] ,
    \top_I.branch[6].l_um_iw[150] ,
    \top_I.branch[6].l_um_iw[149] ,
    \top_I.branch[6].l_um_iw[148] ,
    \top_I.branch[6].l_um_iw[147] ,
    \top_I.branch[6].l_um_iw[146] ,
    \top_I.branch[6].l_um_iw[145] ,
    \top_I.branch[6].l_um_iw[144] ,
    \top_I.branch[6].l_um_iw[143] ,
    \top_I.branch[6].l_um_iw[142] ,
    \top_I.branch[6].l_um_iw[141] ,
    \top_I.branch[6].l_um_iw[140] ,
    \top_I.branch[6].l_um_iw[139] ,
    \top_I.branch[6].l_um_iw[138] ,
    \top_I.branch[6].l_um_iw[137] ,
    \top_I.branch[6].l_um_iw[136] ,
    \top_I.branch[6].l_um_iw[135] ,
    \top_I.branch[6].l_um_iw[134] ,
    \top_I.branch[6].l_um_iw[133] ,
    \top_I.branch[6].l_um_iw[132] ,
    \top_I.branch[6].l_um_iw[131] ,
    \top_I.branch[6].l_um_iw[130] ,
    \top_I.branch[6].l_um_iw[129] ,
    \top_I.branch[6].l_um_iw[128] ,
    \top_I.branch[6].l_um_iw[127] ,
    \top_I.branch[6].l_um_iw[126] ,
    \top_I.branch[6].l_um_iw[125] ,
    \top_I.branch[6].l_um_iw[124] ,
    \top_I.branch[6].l_um_iw[123] ,
    \top_I.branch[6].l_um_iw[122] ,
    \top_I.branch[6].l_um_iw[121] ,
    \top_I.branch[6].l_um_iw[120] ,
    \top_I.branch[6].l_um_iw[119] ,
    \top_I.branch[6].l_um_iw[118] ,
    \top_I.branch[6].l_um_iw[117] ,
    \top_I.branch[6].l_um_iw[116] ,
    \top_I.branch[6].l_um_iw[115] ,
    \top_I.branch[6].l_um_iw[114] ,
    \top_I.branch[6].l_um_iw[113] ,
    \top_I.branch[6].l_um_iw[112] ,
    \top_I.branch[6].l_um_iw[111] ,
    \top_I.branch[6].l_um_iw[110] ,
    \top_I.branch[6].l_um_iw[109] ,
    \top_I.branch[6].l_um_iw[108] ,
    \top_I.branch[6].l_um_iw[107] ,
    \top_I.branch[6].l_um_iw[106] ,
    \top_I.branch[6].l_um_iw[105] ,
    \top_I.branch[6].l_um_iw[104] ,
    \top_I.branch[6].l_um_iw[103] ,
    \top_I.branch[6].l_um_iw[102] ,
    \top_I.branch[6].l_um_iw[101] ,
    \top_I.branch[6].l_um_iw[100] ,
    \top_I.branch[6].l_um_iw[99] ,
    \top_I.branch[6].l_um_iw[98] ,
    \top_I.branch[6].l_um_iw[97] ,
    \top_I.branch[6].l_um_iw[96] ,
    \top_I.branch[6].l_um_iw[95] ,
    \top_I.branch[6].l_um_iw[94] ,
    \top_I.branch[6].l_um_iw[93] ,
    \top_I.branch[6].l_um_iw[92] ,
    \top_I.branch[6].l_um_iw[91] ,
    \top_I.branch[6].l_um_iw[90] ,
    \top_I.branch[6].l_um_iw[89] ,
    \top_I.branch[6].l_um_iw[88] ,
    \top_I.branch[6].l_um_iw[87] ,
    \top_I.branch[6].l_um_iw[86] ,
    \top_I.branch[6].l_um_iw[85] ,
    \top_I.branch[6].l_um_iw[84] ,
    \top_I.branch[6].l_um_iw[83] ,
    \top_I.branch[6].l_um_iw[82] ,
    \top_I.branch[6].l_um_iw[81] ,
    \top_I.branch[6].l_um_iw[80] ,
    \top_I.branch[6].l_um_iw[79] ,
    \top_I.branch[6].l_um_iw[78] ,
    \top_I.branch[6].l_um_iw[77] ,
    \top_I.branch[6].l_um_iw[76] ,
    \top_I.branch[6].l_um_iw[75] ,
    \top_I.branch[6].l_um_iw[74] ,
    \top_I.branch[6].l_um_iw[73] ,
    \top_I.branch[6].l_um_iw[72] ,
    \top_I.branch[6].l_um_iw[71] ,
    \top_I.branch[6].l_um_iw[70] ,
    \top_I.branch[6].l_um_iw[69] ,
    \top_I.branch[6].l_um_iw[68] ,
    \top_I.branch[6].l_um_iw[67] ,
    \top_I.branch[6].l_um_iw[66] ,
    \top_I.branch[6].l_um_iw[65] ,
    \top_I.branch[6].l_um_iw[64] ,
    \top_I.branch[6].l_um_iw[63] ,
    \top_I.branch[6].l_um_iw[62] ,
    \top_I.branch[6].l_um_iw[61] ,
    \top_I.branch[6].l_um_iw[60] ,
    \top_I.branch[6].l_um_iw[59] ,
    \top_I.branch[6].l_um_iw[58] ,
    \top_I.branch[6].l_um_iw[57] ,
    \top_I.branch[6].l_um_iw[56] ,
    \top_I.branch[6].l_um_iw[55] ,
    \top_I.branch[6].l_um_iw[54] ,
    \top_I.branch[6].l_um_iw[53] ,
    \top_I.branch[6].l_um_iw[52] ,
    \top_I.branch[6].l_um_iw[51] ,
    \top_I.branch[6].l_um_iw[50] ,
    \top_I.branch[6].l_um_iw[49] ,
    \top_I.branch[6].l_um_iw[48] ,
    \top_I.branch[6].l_um_iw[47] ,
    \top_I.branch[6].l_um_iw[46] ,
    \top_I.branch[6].l_um_iw[45] ,
    \top_I.branch[6].l_um_iw[44] ,
    \top_I.branch[6].l_um_iw[43] ,
    \top_I.branch[6].l_um_iw[42] ,
    \top_I.branch[6].l_um_iw[41] ,
    \top_I.branch[6].l_um_iw[40] ,
    \top_I.branch[6].l_um_iw[39] ,
    \top_I.branch[6].l_um_iw[38] ,
    \top_I.branch[6].l_um_iw[37] ,
    \top_I.branch[6].l_um_iw[36] ,
    \top_I.branch[6].l_um_iw[35] ,
    \top_I.branch[6].l_um_iw[34] ,
    \top_I.branch[6].l_um_iw[33] ,
    \top_I.branch[6].l_um_iw[32] ,
    \top_I.branch[6].l_um_iw[31] ,
    \top_I.branch[6].l_um_iw[30] ,
    \top_I.branch[6].l_um_iw[29] ,
    \top_I.branch[6].l_um_iw[28] ,
    \top_I.branch[6].l_um_iw[27] ,
    \top_I.branch[6].l_um_iw[26] ,
    \top_I.branch[6].l_um_iw[25] ,
    \top_I.branch[6].l_um_iw[24] ,
    \top_I.branch[6].l_um_iw[23] ,
    \top_I.branch[6].l_um_iw[22] ,
    \top_I.branch[6].l_um_iw[21] ,
    \top_I.branch[6].l_um_iw[20] ,
    \top_I.branch[6].l_um_iw[19] ,
    \top_I.branch[6].l_um_iw[18] ,
    \top_I.branch[6].l_um_iw[17] ,
    \top_I.branch[6].l_um_iw[16] ,
    \top_I.branch[6].l_um_iw[15] ,
    \top_I.branch[6].l_um_iw[14] ,
    \top_I.branch[6].l_um_iw[13] ,
    \top_I.branch[6].l_um_iw[12] ,
    \top_I.branch[6].l_um_iw[11] ,
    \top_I.branch[6].l_um_iw[10] ,
    \top_I.branch[6].l_um_iw[9] ,
    \top_I.branch[6].l_um_iw[8] ,
    \top_I.branch[6].l_um_iw[7] ,
    \top_I.branch[6].l_um_iw[6] ,
    \top_I.branch[6].l_um_iw[5] ,
    \top_I.branch[6].l_um_iw[4] ,
    \top_I.branch[6].l_um_iw[3] ,
    \top_I.branch[6].l_um_iw[2] ,
    \top_I.branch[6].l_um_iw[1] ,
    \top_I.branch[6].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[1] ,
    \top_I.branch[6].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[15] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[14] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[13] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[12] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[11] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[10] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[9] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[8] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[7] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[6] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[5] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[4] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[3] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].l_um_k_zero[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[6].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] ,
    \top_I.branch[6].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[7].col_um[0].um_top_I.block_7_16.tt_um_I  (.clk(\top_I.branch[7].l_um_iw[18] ),
    .ena(\top_I.branch[7].l_um_ena[1] ),
    .rst_n(\top_I.branch[7].l_um_iw[19] ),
    .ui_in({\top_I.branch[7].l_um_iw[27] ,
    \top_I.branch[7].l_um_iw[26] ,
    \top_I.branch[7].l_um_iw[25] ,
    \top_I.branch[7].l_um_iw[24] ,
    \top_I.branch[7].l_um_iw[23] ,
    \top_I.branch[7].l_um_iw[22] ,
    \top_I.branch[7].l_um_iw[21] ,
    \top_I.branch[7].l_um_iw[20] }),
    .uio_in({\top_I.branch[7].l_um_iw[35] ,
    \top_I.branch[7].l_um_iw[34] ,
    \top_I.branch[7].l_um_iw[33] ,
    \top_I.branch[7].l_um_iw[32] ,
    \top_I.branch[7].l_um_iw[31] ,
    \top_I.branch[7].l_um_iw[30] ,
    \top_I.branch[7].l_um_iw[29] ,
    \top_I.branch[7].l_um_iw[28] }),
    .uio_oe({\top_I.branch[7].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[0] }),
    .uio_out({\top_I.branch[7].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[0] }),
    .uo_out({\top_I.branch[7].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[0] }));
 tt_mux \top_I.branch[7].mux_I  (.k_one(\top_I.branch[7].l_k_one ),
    .k_zero(\top_I.branch[7].l_k_zero ),
    .addr({\top_I.branch[7].l_k_zero ,
    \top_I.branch[7].l_k_zero ,
    \top_I.branch[7].l_k_one ,
    \top_I.branch[7].l_k_one ,
    \top_I.branch[7].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[7].l_um_ena[15] ,
    \top_I.branch[7].l_um_ena[14] ,
    \top_I.branch[7].l_um_ena[13] ,
    \top_I.branch[7].l_um_ena[12] ,
    \top_I.branch[7].l_um_ena[11] ,
    \top_I.branch[7].l_um_ena[10] ,
    \top_I.branch[7].l_um_ena[9] ,
    \top_I.branch[7].l_um_ena[8] ,
    \top_I.branch[7].l_um_ena[7] ,
    \top_I.branch[7].l_um_ena[6] ,
    \top_I.branch[7].l_um_ena[5] ,
    \top_I.branch[7].l_um_ena[4] ,
    \top_I.branch[7].l_um_ena[3] ,
    \top_I.branch[7].l_um_ena[2] ,
    \top_I.branch[7].l_um_ena[1] ,
    \top_I.branch[7].l_um_ena[0] }),
    .um_iw({\top_I.branch[7].l_um_iw[287] ,
    \top_I.branch[7].l_um_iw[286] ,
    \top_I.branch[7].l_um_iw[285] ,
    \top_I.branch[7].l_um_iw[284] ,
    \top_I.branch[7].l_um_iw[283] ,
    \top_I.branch[7].l_um_iw[282] ,
    \top_I.branch[7].l_um_iw[281] ,
    \top_I.branch[7].l_um_iw[280] ,
    \top_I.branch[7].l_um_iw[279] ,
    \top_I.branch[7].l_um_iw[278] ,
    \top_I.branch[7].l_um_iw[277] ,
    \top_I.branch[7].l_um_iw[276] ,
    \top_I.branch[7].l_um_iw[275] ,
    \top_I.branch[7].l_um_iw[274] ,
    \top_I.branch[7].l_um_iw[273] ,
    \top_I.branch[7].l_um_iw[272] ,
    \top_I.branch[7].l_um_iw[271] ,
    \top_I.branch[7].l_um_iw[270] ,
    \top_I.branch[7].l_um_iw[269] ,
    \top_I.branch[7].l_um_iw[268] ,
    \top_I.branch[7].l_um_iw[267] ,
    \top_I.branch[7].l_um_iw[266] ,
    \top_I.branch[7].l_um_iw[265] ,
    \top_I.branch[7].l_um_iw[264] ,
    \top_I.branch[7].l_um_iw[263] ,
    \top_I.branch[7].l_um_iw[262] ,
    \top_I.branch[7].l_um_iw[261] ,
    \top_I.branch[7].l_um_iw[260] ,
    \top_I.branch[7].l_um_iw[259] ,
    \top_I.branch[7].l_um_iw[258] ,
    \top_I.branch[7].l_um_iw[257] ,
    \top_I.branch[7].l_um_iw[256] ,
    \top_I.branch[7].l_um_iw[255] ,
    \top_I.branch[7].l_um_iw[254] ,
    \top_I.branch[7].l_um_iw[253] ,
    \top_I.branch[7].l_um_iw[252] ,
    \top_I.branch[7].l_um_iw[251] ,
    \top_I.branch[7].l_um_iw[250] ,
    \top_I.branch[7].l_um_iw[249] ,
    \top_I.branch[7].l_um_iw[248] ,
    \top_I.branch[7].l_um_iw[247] ,
    \top_I.branch[7].l_um_iw[246] ,
    \top_I.branch[7].l_um_iw[245] ,
    \top_I.branch[7].l_um_iw[244] ,
    \top_I.branch[7].l_um_iw[243] ,
    \top_I.branch[7].l_um_iw[242] ,
    \top_I.branch[7].l_um_iw[241] ,
    \top_I.branch[7].l_um_iw[240] ,
    \top_I.branch[7].l_um_iw[239] ,
    \top_I.branch[7].l_um_iw[238] ,
    \top_I.branch[7].l_um_iw[237] ,
    \top_I.branch[7].l_um_iw[236] ,
    \top_I.branch[7].l_um_iw[235] ,
    \top_I.branch[7].l_um_iw[234] ,
    \top_I.branch[7].l_um_iw[233] ,
    \top_I.branch[7].l_um_iw[232] ,
    \top_I.branch[7].l_um_iw[231] ,
    \top_I.branch[7].l_um_iw[230] ,
    \top_I.branch[7].l_um_iw[229] ,
    \top_I.branch[7].l_um_iw[228] ,
    \top_I.branch[7].l_um_iw[227] ,
    \top_I.branch[7].l_um_iw[226] ,
    \top_I.branch[7].l_um_iw[225] ,
    \top_I.branch[7].l_um_iw[224] ,
    \top_I.branch[7].l_um_iw[223] ,
    \top_I.branch[7].l_um_iw[222] ,
    \top_I.branch[7].l_um_iw[221] ,
    \top_I.branch[7].l_um_iw[220] ,
    \top_I.branch[7].l_um_iw[219] ,
    \top_I.branch[7].l_um_iw[218] ,
    \top_I.branch[7].l_um_iw[217] ,
    \top_I.branch[7].l_um_iw[216] ,
    \top_I.branch[7].l_um_iw[215] ,
    \top_I.branch[7].l_um_iw[214] ,
    \top_I.branch[7].l_um_iw[213] ,
    \top_I.branch[7].l_um_iw[212] ,
    \top_I.branch[7].l_um_iw[211] ,
    \top_I.branch[7].l_um_iw[210] ,
    \top_I.branch[7].l_um_iw[209] ,
    \top_I.branch[7].l_um_iw[208] ,
    \top_I.branch[7].l_um_iw[207] ,
    \top_I.branch[7].l_um_iw[206] ,
    \top_I.branch[7].l_um_iw[205] ,
    \top_I.branch[7].l_um_iw[204] ,
    \top_I.branch[7].l_um_iw[203] ,
    \top_I.branch[7].l_um_iw[202] ,
    \top_I.branch[7].l_um_iw[201] ,
    \top_I.branch[7].l_um_iw[200] ,
    \top_I.branch[7].l_um_iw[199] ,
    \top_I.branch[7].l_um_iw[198] ,
    \top_I.branch[7].l_um_iw[197] ,
    \top_I.branch[7].l_um_iw[196] ,
    \top_I.branch[7].l_um_iw[195] ,
    \top_I.branch[7].l_um_iw[194] ,
    \top_I.branch[7].l_um_iw[193] ,
    \top_I.branch[7].l_um_iw[192] ,
    \top_I.branch[7].l_um_iw[191] ,
    \top_I.branch[7].l_um_iw[190] ,
    \top_I.branch[7].l_um_iw[189] ,
    \top_I.branch[7].l_um_iw[188] ,
    \top_I.branch[7].l_um_iw[187] ,
    \top_I.branch[7].l_um_iw[186] ,
    \top_I.branch[7].l_um_iw[185] ,
    \top_I.branch[7].l_um_iw[184] ,
    \top_I.branch[7].l_um_iw[183] ,
    \top_I.branch[7].l_um_iw[182] ,
    \top_I.branch[7].l_um_iw[181] ,
    \top_I.branch[7].l_um_iw[180] ,
    \top_I.branch[7].l_um_iw[179] ,
    \top_I.branch[7].l_um_iw[178] ,
    \top_I.branch[7].l_um_iw[177] ,
    \top_I.branch[7].l_um_iw[176] ,
    \top_I.branch[7].l_um_iw[175] ,
    \top_I.branch[7].l_um_iw[174] ,
    \top_I.branch[7].l_um_iw[173] ,
    \top_I.branch[7].l_um_iw[172] ,
    \top_I.branch[7].l_um_iw[171] ,
    \top_I.branch[7].l_um_iw[170] ,
    \top_I.branch[7].l_um_iw[169] ,
    \top_I.branch[7].l_um_iw[168] ,
    \top_I.branch[7].l_um_iw[167] ,
    \top_I.branch[7].l_um_iw[166] ,
    \top_I.branch[7].l_um_iw[165] ,
    \top_I.branch[7].l_um_iw[164] ,
    \top_I.branch[7].l_um_iw[163] ,
    \top_I.branch[7].l_um_iw[162] ,
    \top_I.branch[7].l_um_iw[161] ,
    \top_I.branch[7].l_um_iw[160] ,
    \top_I.branch[7].l_um_iw[159] ,
    \top_I.branch[7].l_um_iw[158] ,
    \top_I.branch[7].l_um_iw[157] ,
    \top_I.branch[7].l_um_iw[156] ,
    \top_I.branch[7].l_um_iw[155] ,
    \top_I.branch[7].l_um_iw[154] ,
    \top_I.branch[7].l_um_iw[153] ,
    \top_I.branch[7].l_um_iw[152] ,
    \top_I.branch[7].l_um_iw[151] ,
    \top_I.branch[7].l_um_iw[150] ,
    \top_I.branch[7].l_um_iw[149] ,
    \top_I.branch[7].l_um_iw[148] ,
    \top_I.branch[7].l_um_iw[147] ,
    \top_I.branch[7].l_um_iw[146] ,
    \top_I.branch[7].l_um_iw[145] ,
    \top_I.branch[7].l_um_iw[144] ,
    \top_I.branch[7].l_um_iw[143] ,
    \top_I.branch[7].l_um_iw[142] ,
    \top_I.branch[7].l_um_iw[141] ,
    \top_I.branch[7].l_um_iw[140] ,
    \top_I.branch[7].l_um_iw[139] ,
    \top_I.branch[7].l_um_iw[138] ,
    \top_I.branch[7].l_um_iw[137] ,
    \top_I.branch[7].l_um_iw[136] ,
    \top_I.branch[7].l_um_iw[135] ,
    \top_I.branch[7].l_um_iw[134] ,
    \top_I.branch[7].l_um_iw[133] ,
    \top_I.branch[7].l_um_iw[132] ,
    \top_I.branch[7].l_um_iw[131] ,
    \top_I.branch[7].l_um_iw[130] ,
    \top_I.branch[7].l_um_iw[129] ,
    \top_I.branch[7].l_um_iw[128] ,
    \top_I.branch[7].l_um_iw[127] ,
    \top_I.branch[7].l_um_iw[126] ,
    \top_I.branch[7].l_um_iw[125] ,
    \top_I.branch[7].l_um_iw[124] ,
    \top_I.branch[7].l_um_iw[123] ,
    \top_I.branch[7].l_um_iw[122] ,
    \top_I.branch[7].l_um_iw[121] ,
    \top_I.branch[7].l_um_iw[120] ,
    \top_I.branch[7].l_um_iw[119] ,
    \top_I.branch[7].l_um_iw[118] ,
    \top_I.branch[7].l_um_iw[117] ,
    \top_I.branch[7].l_um_iw[116] ,
    \top_I.branch[7].l_um_iw[115] ,
    \top_I.branch[7].l_um_iw[114] ,
    \top_I.branch[7].l_um_iw[113] ,
    \top_I.branch[7].l_um_iw[112] ,
    \top_I.branch[7].l_um_iw[111] ,
    \top_I.branch[7].l_um_iw[110] ,
    \top_I.branch[7].l_um_iw[109] ,
    \top_I.branch[7].l_um_iw[108] ,
    \top_I.branch[7].l_um_iw[107] ,
    \top_I.branch[7].l_um_iw[106] ,
    \top_I.branch[7].l_um_iw[105] ,
    \top_I.branch[7].l_um_iw[104] ,
    \top_I.branch[7].l_um_iw[103] ,
    \top_I.branch[7].l_um_iw[102] ,
    \top_I.branch[7].l_um_iw[101] ,
    \top_I.branch[7].l_um_iw[100] ,
    \top_I.branch[7].l_um_iw[99] ,
    \top_I.branch[7].l_um_iw[98] ,
    \top_I.branch[7].l_um_iw[97] ,
    \top_I.branch[7].l_um_iw[96] ,
    \top_I.branch[7].l_um_iw[95] ,
    \top_I.branch[7].l_um_iw[94] ,
    \top_I.branch[7].l_um_iw[93] ,
    \top_I.branch[7].l_um_iw[92] ,
    \top_I.branch[7].l_um_iw[91] ,
    \top_I.branch[7].l_um_iw[90] ,
    \top_I.branch[7].l_um_iw[89] ,
    \top_I.branch[7].l_um_iw[88] ,
    \top_I.branch[7].l_um_iw[87] ,
    \top_I.branch[7].l_um_iw[86] ,
    \top_I.branch[7].l_um_iw[85] ,
    \top_I.branch[7].l_um_iw[84] ,
    \top_I.branch[7].l_um_iw[83] ,
    \top_I.branch[7].l_um_iw[82] ,
    \top_I.branch[7].l_um_iw[81] ,
    \top_I.branch[7].l_um_iw[80] ,
    \top_I.branch[7].l_um_iw[79] ,
    \top_I.branch[7].l_um_iw[78] ,
    \top_I.branch[7].l_um_iw[77] ,
    \top_I.branch[7].l_um_iw[76] ,
    \top_I.branch[7].l_um_iw[75] ,
    \top_I.branch[7].l_um_iw[74] ,
    \top_I.branch[7].l_um_iw[73] ,
    \top_I.branch[7].l_um_iw[72] ,
    \top_I.branch[7].l_um_iw[71] ,
    \top_I.branch[7].l_um_iw[70] ,
    \top_I.branch[7].l_um_iw[69] ,
    \top_I.branch[7].l_um_iw[68] ,
    \top_I.branch[7].l_um_iw[67] ,
    \top_I.branch[7].l_um_iw[66] ,
    \top_I.branch[7].l_um_iw[65] ,
    \top_I.branch[7].l_um_iw[64] ,
    \top_I.branch[7].l_um_iw[63] ,
    \top_I.branch[7].l_um_iw[62] ,
    \top_I.branch[7].l_um_iw[61] ,
    \top_I.branch[7].l_um_iw[60] ,
    \top_I.branch[7].l_um_iw[59] ,
    \top_I.branch[7].l_um_iw[58] ,
    \top_I.branch[7].l_um_iw[57] ,
    \top_I.branch[7].l_um_iw[56] ,
    \top_I.branch[7].l_um_iw[55] ,
    \top_I.branch[7].l_um_iw[54] ,
    \top_I.branch[7].l_um_iw[53] ,
    \top_I.branch[7].l_um_iw[52] ,
    \top_I.branch[7].l_um_iw[51] ,
    \top_I.branch[7].l_um_iw[50] ,
    \top_I.branch[7].l_um_iw[49] ,
    \top_I.branch[7].l_um_iw[48] ,
    \top_I.branch[7].l_um_iw[47] ,
    \top_I.branch[7].l_um_iw[46] ,
    \top_I.branch[7].l_um_iw[45] ,
    \top_I.branch[7].l_um_iw[44] ,
    \top_I.branch[7].l_um_iw[43] ,
    \top_I.branch[7].l_um_iw[42] ,
    \top_I.branch[7].l_um_iw[41] ,
    \top_I.branch[7].l_um_iw[40] ,
    \top_I.branch[7].l_um_iw[39] ,
    \top_I.branch[7].l_um_iw[38] ,
    \top_I.branch[7].l_um_iw[37] ,
    \top_I.branch[7].l_um_iw[36] ,
    \top_I.branch[7].l_um_iw[35] ,
    \top_I.branch[7].l_um_iw[34] ,
    \top_I.branch[7].l_um_iw[33] ,
    \top_I.branch[7].l_um_iw[32] ,
    \top_I.branch[7].l_um_iw[31] ,
    \top_I.branch[7].l_um_iw[30] ,
    \top_I.branch[7].l_um_iw[29] ,
    \top_I.branch[7].l_um_iw[28] ,
    \top_I.branch[7].l_um_iw[27] ,
    \top_I.branch[7].l_um_iw[26] ,
    \top_I.branch[7].l_um_iw[25] ,
    \top_I.branch[7].l_um_iw[24] ,
    \top_I.branch[7].l_um_iw[23] ,
    \top_I.branch[7].l_um_iw[22] ,
    \top_I.branch[7].l_um_iw[21] ,
    \top_I.branch[7].l_um_iw[20] ,
    \top_I.branch[7].l_um_iw[19] ,
    \top_I.branch[7].l_um_iw[18] ,
    \top_I.branch[7].l_um_iw[17] ,
    \top_I.branch[7].l_um_iw[16] ,
    \top_I.branch[7].l_um_iw[15] ,
    \top_I.branch[7].l_um_iw[14] ,
    \top_I.branch[7].l_um_iw[13] ,
    \top_I.branch[7].l_um_iw[12] ,
    \top_I.branch[7].l_um_iw[11] ,
    \top_I.branch[7].l_um_iw[10] ,
    \top_I.branch[7].l_um_iw[9] ,
    \top_I.branch[7].l_um_iw[8] ,
    \top_I.branch[7].l_um_iw[7] ,
    \top_I.branch[7].l_um_iw[6] ,
    \top_I.branch[7].l_um_iw[5] ,
    \top_I.branch[7].l_um_iw[4] ,
    \top_I.branch[7].l_um_iw[3] ,
    \top_I.branch[7].l_um_iw[2] ,
    \top_I.branch[7].l_um_iw[1] ,
    \top_I.branch[7].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[1] ,
    \top_I.branch[7].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[15] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[14] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[13] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[12] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[11] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[10] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[9] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[8] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[7] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[6] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[5] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[4] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[3] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].l_um_k_zero[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_oe[0] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uio_out[0] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[7] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[6] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[5] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[4] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[3] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[2] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[1] ,
    \top_I.branch[7].col_um[0].um_top_I.uo_out[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] ,
    \top_I.branch[7].l_um_k_zero[0] }));
 tt_um_loopback \top_I.branch[8].col_um[0].um_bot_I.block_8_0.tt_um_I  (.clk(\top_I.branch[8].l_um_iw[0] ),
    .ena(\top_I.branch[8].l_um_ena[0] ),
    .rst_n(\top_I.branch[8].l_um_iw[1] ),
    .ui_in({\top_I.branch[8].l_um_iw[9] ,
    \top_I.branch[8].l_um_iw[8] ,
    \top_I.branch[8].l_um_iw[7] ,
    \top_I.branch[8].l_um_iw[6] ,
    \top_I.branch[8].l_um_iw[5] ,
    \top_I.branch[8].l_um_iw[4] ,
    \top_I.branch[8].l_um_iw[3] ,
    \top_I.branch[8].l_um_iw[2] }),
    .uio_in({\top_I.branch[8].l_um_iw[17] ,
    \top_I.branch[8].l_um_iw[16] ,
    \top_I.branch[8].l_um_iw[15] ,
    \top_I.branch[8].l_um_iw[14] ,
    \top_I.branch[8].l_um_iw[13] ,
    \top_I.branch[8].l_um_iw[12] ,
    \top_I.branch[8].l_um_iw[11] ,
    \top_I.branch[8].l_um_iw[10] }),
    .uio_oe({\top_I.branch[8].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[8].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[8].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[8].mux_I  (.k_one(\top_I.branch[8].l_k_one ),
    .k_zero(\top_I.branch[8].l_k_zero ),
    .addr({\top_I.branch[8].l_k_zero ,
    \top_I.branch[8].l_k_one ,
    \top_I.branch[8].l_k_zero ,
    \top_I.branch[8].l_k_zero ,
    \top_I.branch[8].l_k_zero }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[8].l_um_ena[15] ,
    \top_I.branch[8].l_um_ena[14] ,
    \top_I.branch[8].l_um_ena[13] ,
    \top_I.branch[8].l_um_ena[12] ,
    \top_I.branch[8].l_um_ena[11] ,
    \top_I.branch[8].l_um_ena[10] ,
    \top_I.branch[8].l_um_ena[9] ,
    \top_I.branch[8].l_um_ena[8] ,
    \top_I.branch[8].l_um_ena[7] ,
    \top_I.branch[8].l_um_ena[6] ,
    \top_I.branch[8].l_um_ena[5] ,
    \top_I.branch[8].l_um_ena[4] ,
    \top_I.branch[8].l_um_ena[3] ,
    \top_I.branch[8].l_um_ena[2] ,
    \top_I.branch[8].l_um_ena[1] ,
    \top_I.branch[8].l_um_ena[0] }),
    .um_iw({\top_I.branch[8].l_um_iw[287] ,
    \top_I.branch[8].l_um_iw[286] ,
    \top_I.branch[8].l_um_iw[285] ,
    \top_I.branch[8].l_um_iw[284] ,
    \top_I.branch[8].l_um_iw[283] ,
    \top_I.branch[8].l_um_iw[282] ,
    \top_I.branch[8].l_um_iw[281] ,
    \top_I.branch[8].l_um_iw[280] ,
    \top_I.branch[8].l_um_iw[279] ,
    \top_I.branch[8].l_um_iw[278] ,
    \top_I.branch[8].l_um_iw[277] ,
    \top_I.branch[8].l_um_iw[276] ,
    \top_I.branch[8].l_um_iw[275] ,
    \top_I.branch[8].l_um_iw[274] ,
    \top_I.branch[8].l_um_iw[273] ,
    \top_I.branch[8].l_um_iw[272] ,
    \top_I.branch[8].l_um_iw[271] ,
    \top_I.branch[8].l_um_iw[270] ,
    \top_I.branch[8].l_um_iw[269] ,
    \top_I.branch[8].l_um_iw[268] ,
    \top_I.branch[8].l_um_iw[267] ,
    \top_I.branch[8].l_um_iw[266] ,
    \top_I.branch[8].l_um_iw[265] ,
    \top_I.branch[8].l_um_iw[264] ,
    \top_I.branch[8].l_um_iw[263] ,
    \top_I.branch[8].l_um_iw[262] ,
    \top_I.branch[8].l_um_iw[261] ,
    \top_I.branch[8].l_um_iw[260] ,
    \top_I.branch[8].l_um_iw[259] ,
    \top_I.branch[8].l_um_iw[258] ,
    \top_I.branch[8].l_um_iw[257] ,
    \top_I.branch[8].l_um_iw[256] ,
    \top_I.branch[8].l_um_iw[255] ,
    \top_I.branch[8].l_um_iw[254] ,
    \top_I.branch[8].l_um_iw[253] ,
    \top_I.branch[8].l_um_iw[252] ,
    \top_I.branch[8].l_um_iw[251] ,
    \top_I.branch[8].l_um_iw[250] ,
    \top_I.branch[8].l_um_iw[249] ,
    \top_I.branch[8].l_um_iw[248] ,
    \top_I.branch[8].l_um_iw[247] ,
    \top_I.branch[8].l_um_iw[246] ,
    \top_I.branch[8].l_um_iw[245] ,
    \top_I.branch[8].l_um_iw[244] ,
    \top_I.branch[8].l_um_iw[243] ,
    \top_I.branch[8].l_um_iw[242] ,
    \top_I.branch[8].l_um_iw[241] ,
    \top_I.branch[8].l_um_iw[240] ,
    \top_I.branch[8].l_um_iw[239] ,
    \top_I.branch[8].l_um_iw[238] ,
    \top_I.branch[8].l_um_iw[237] ,
    \top_I.branch[8].l_um_iw[236] ,
    \top_I.branch[8].l_um_iw[235] ,
    \top_I.branch[8].l_um_iw[234] ,
    \top_I.branch[8].l_um_iw[233] ,
    \top_I.branch[8].l_um_iw[232] ,
    \top_I.branch[8].l_um_iw[231] ,
    \top_I.branch[8].l_um_iw[230] ,
    \top_I.branch[8].l_um_iw[229] ,
    \top_I.branch[8].l_um_iw[228] ,
    \top_I.branch[8].l_um_iw[227] ,
    \top_I.branch[8].l_um_iw[226] ,
    \top_I.branch[8].l_um_iw[225] ,
    \top_I.branch[8].l_um_iw[224] ,
    \top_I.branch[8].l_um_iw[223] ,
    \top_I.branch[8].l_um_iw[222] ,
    \top_I.branch[8].l_um_iw[221] ,
    \top_I.branch[8].l_um_iw[220] ,
    \top_I.branch[8].l_um_iw[219] ,
    \top_I.branch[8].l_um_iw[218] ,
    \top_I.branch[8].l_um_iw[217] ,
    \top_I.branch[8].l_um_iw[216] ,
    \top_I.branch[8].l_um_iw[215] ,
    \top_I.branch[8].l_um_iw[214] ,
    \top_I.branch[8].l_um_iw[213] ,
    \top_I.branch[8].l_um_iw[212] ,
    \top_I.branch[8].l_um_iw[211] ,
    \top_I.branch[8].l_um_iw[210] ,
    \top_I.branch[8].l_um_iw[209] ,
    \top_I.branch[8].l_um_iw[208] ,
    \top_I.branch[8].l_um_iw[207] ,
    \top_I.branch[8].l_um_iw[206] ,
    \top_I.branch[8].l_um_iw[205] ,
    \top_I.branch[8].l_um_iw[204] ,
    \top_I.branch[8].l_um_iw[203] ,
    \top_I.branch[8].l_um_iw[202] ,
    \top_I.branch[8].l_um_iw[201] ,
    \top_I.branch[8].l_um_iw[200] ,
    \top_I.branch[8].l_um_iw[199] ,
    \top_I.branch[8].l_um_iw[198] ,
    \top_I.branch[8].l_um_iw[197] ,
    \top_I.branch[8].l_um_iw[196] ,
    \top_I.branch[8].l_um_iw[195] ,
    \top_I.branch[8].l_um_iw[194] ,
    \top_I.branch[8].l_um_iw[193] ,
    \top_I.branch[8].l_um_iw[192] ,
    \top_I.branch[8].l_um_iw[191] ,
    \top_I.branch[8].l_um_iw[190] ,
    \top_I.branch[8].l_um_iw[189] ,
    \top_I.branch[8].l_um_iw[188] ,
    \top_I.branch[8].l_um_iw[187] ,
    \top_I.branch[8].l_um_iw[186] ,
    \top_I.branch[8].l_um_iw[185] ,
    \top_I.branch[8].l_um_iw[184] ,
    \top_I.branch[8].l_um_iw[183] ,
    \top_I.branch[8].l_um_iw[182] ,
    \top_I.branch[8].l_um_iw[181] ,
    \top_I.branch[8].l_um_iw[180] ,
    \top_I.branch[8].l_um_iw[179] ,
    \top_I.branch[8].l_um_iw[178] ,
    \top_I.branch[8].l_um_iw[177] ,
    \top_I.branch[8].l_um_iw[176] ,
    \top_I.branch[8].l_um_iw[175] ,
    \top_I.branch[8].l_um_iw[174] ,
    \top_I.branch[8].l_um_iw[173] ,
    \top_I.branch[8].l_um_iw[172] ,
    \top_I.branch[8].l_um_iw[171] ,
    \top_I.branch[8].l_um_iw[170] ,
    \top_I.branch[8].l_um_iw[169] ,
    \top_I.branch[8].l_um_iw[168] ,
    \top_I.branch[8].l_um_iw[167] ,
    \top_I.branch[8].l_um_iw[166] ,
    \top_I.branch[8].l_um_iw[165] ,
    \top_I.branch[8].l_um_iw[164] ,
    \top_I.branch[8].l_um_iw[163] ,
    \top_I.branch[8].l_um_iw[162] ,
    \top_I.branch[8].l_um_iw[161] ,
    \top_I.branch[8].l_um_iw[160] ,
    \top_I.branch[8].l_um_iw[159] ,
    \top_I.branch[8].l_um_iw[158] ,
    \top_I.branch[8].l_um_iw[157] ,
    \top_I.branch[8].l_um_iw[156] ,
    \top_I.branch[8].l_um_iw[155] ,
    \top_I.branch[8].l_um_iw[154] ,
    \top_I.branch[8].l_um_iw[153] ,
    \top_I.branch[8].l_um_iw[152] ,
    \top_I.branch[8].l_um_iw[151] ,
    \top_I.branch[8].l_um_iw[150] ,
    \top_I.branch[8].l_um_iw[149] ,
    \top_I.branch[8].l_um_iw[148] ,
    \top_I.branch[8].l_um_iw[147] ,
    \top_I.branch[8].l_um_iw[146] ,
    \top_I.branch[8].l_um_iw[145] ,
    \top_I.branch[8].l_um_iw[144] ,
    \top_I.branch[8].l_um_iw[143] ,
    \top_I.branch[8].l_um_iw[142] ,
    \top_I.branch[8].l_um_iw[141] ,
    \top_I.branch[8].l_um_iw[140] ,
    \top_I.branch[8].l_um_iw[139] ,
    \top_I.branch[8].l_um_iw[138] ,
    \top_I.branch[8].l_um_iw[137] ,
    \top_I.branch[8].l_um_iw[136] ,
    \top_I.branch[8].l_um_iw[135] ,
    \top_I.branch[8].l_um_iw[134] ,
    \top_I.branch[8].l_um_iw[133] ,
    \top_I.branch[8].l_um_iw[132] ,
    \top_I.branch[8].l_um_iw[131] ,
    \top_I.branch[8].l_um_iw[130] ,
    \top_I.branch[8].l_um_iw[129] ,
    \top_I.branch[8].l_um_iw[128] ,
    \top_I.branch[8].l_um_iw[127] ,
    \top_I.branch[8].l_um_iw[126] ,
    \top_I.branch[8].l_um_iw[125] ,
    \top_I.branch[8].l_um_iw[124] ,
    \top_I.branch[8].l_um_iw[123] ,
    \top_I.branch[8].l_um_iw[122] ,
    \top_I.branch[8].l_um_iw[121] ,
    \top_I.branch[8].l_um_iw[120] ,
    \top_I.branch[8].l_um_iw[119] ,
    \top_I.branch[8].l_um_iw[118] ,
    \top_I.branch[8].l_um_iw[117] ,
    \top_I.branch[8].l_um_iw[116] ,
    \top_I.branch[8].l_um_iw[115] ,
    \top_I.branch[8].l_um_iw[114] ,
    \top_I.branch[8].l_um_iw[113] ,
    \top_I.branch[8].l_um_iw[112] ,
    \top_I.branch[8].l_um_iw[111] ,
    \top_I.branch[8].l_um_iw[110] ,
    \top_I.branch[8].l_um_iw[109] ,
    \top_I.branch[8].l_um_iw[108] ,
    \top_I.branch[8].l_um_iw[107] ,
    \top_I.branch[8].l_um_iw[106] ,
    \top_I.branch[8].l_um_iw[105] ,
    \top_I.branch[8].l_um_iw[104] ,
    \top_I.branch[8].l_um_iw[103] ,
    \top_I.branch[8].l_um_iw[102] ,
    \top_I.branch[8].l_um_iw[101] ,
    \top_I.branch[8].l_um_iw[100] ,
    \top_I.branch[8].l_um_iw[99] ,
    \top_I.branch[8].l_um_iw[98] ,
    \top_I.branch[8].l_um_iw[97] ,
    \top_I.branch[8].l_um_iw[96] ,
    \top_I.branch[8].l_um_iw[95] ,
    \top_I.branch[8].l_um_iw[94] ,
    \top_I.branch[8].l_um_iw[93] ,
    \top_I.branch[8].l_um_iw[92] ,
    \top_I.branch[8].l_um_iw[91] ,
    \top_I.branch[8].l_um_iw[90] ,
    \top_I.branch[8].l_um_iw[89] ,
    \top_I.branch[8].l_um_iw[88] ,
    \top_I.branch[8].l_um_iw[87] ,
    \top_I.branch[8].l_um_iw[86] ,
    \top_I.branch[8].l_um_iw[85] ,
    \top_I.branch[8].l_um_iw[84] ,
    \top_I.branch[8].l_um_iw[83] ,
    \top_I.branch[8].l_um_iw[82] ,
    \top_I.branch[8].l_um_iw[81] ,
    \top_I.branch[8].l_um_iw[80] ,
    \top_I.branch[8].l_um_iw[79] ,
    \top_I.branch[8].l_um_iw[78] ,
    \top_I.branch[8].l_um_iw[77] ,
    \top_I.branch[8].l_um_iw[76] ,
    \top_I.branch[8].l_um_iw[75] ,
    \top_I.branch[8].l_um_iw[74] ,
    \top_I.branch[8].l_um_iw[73] ,
    \top_I.branch[8].l_um_iw[72] ,
    \top_I.branch[8].l_um_iw[71] ,
    \top_I.branch[8].l_um_iw[70] ,
    \top_I.branch[8].l_um_iw[69] ,
    \top_I.branch[8].l_um_iw[68] ,
    \top_I.branch[8].l_um_iw[67] ,
    \top_I.branch[8].l_um_iw[66] ,
    \top_I.branch[8].l_um_iw[65] ,
    \top_I.branch[8].l_um_iw[64] ,
    \top_I.branch[8].l_um_iw[63] ,
    \top_I.branch[8].l_um_iw[62] ,
    \top_I.branch[8].l_um_iw[61] ,
    \top_I.branch[8].l_um_iw[60] ,
    \top_I.branch[8].l_um_iw[59] ,
    \top_I.branch[8].l_um_iw[58] ,
    \top_I.branch[8].l_um_iw[57] ,
    \top_I.branch[8].l_um_iw[56] ,
    \top_I.branch[8].l_um_iw[55] ,
    \top_I.branch[8].l_um_iw[54] ,
    \top_I.branch[8].l_um_iw[53] ,
    \top_I.branch[8].l_um_iw[52] ,
    \top_I.branch[8].l_um_iw[51] ,
    \top_I.branch[8].l_um_iw[50] ,
    \top_I.branch[8].l_um_iw[49] ,
    \top_I.branch[8].l_um_iw[48] ,
    \top_I.branch[8].l_um_iw[47] ,
    \top_I.branch[8].l_um_iw[46] ,
    \top_I.branch[8].l_um_iw[45] ,
    \top_I.branch[8].l_um_iw[44] ,
    \top_I.branch[8].l_um_iw[43] ,
    \top_I.branch[8].l_um_iw[42] ,
    \top_I.branch[8].l_um_iw[41] ,
    \top_I.branch[8].l_um_iw[40] ,
    \top_I.branch[8].l_um_iw[39] ,
    \top_I.branch[8].l_um_iw[38] ,
    \top_I.branch[8].l_um_iw[37] ,
    \top_I.branch[8].l_um_iw[36] ,
    \top_I.branch[8].l_um_iw[35] ,
    \top_I.branch[8].l_um_iw[34] ,
    \top_I.branch[8].l_um_iw[33] ,
    \top_I.branch[8].l_um_iw[32] ,
    \top_I.branch[8].l_um_iw[31] ,
    \top_I.branch[8].l_um_iw[30] ,
    \top_I.branch[8].l_um_iw[29] ,
    \top_I.branch[8].l_um_iw[28] ,
    \top_I.branch[8].l_um_iw[27] ,
    \top_I.branch[8].l_um_iw[26] ,
    \top_I.branch[8].l_um_iw[25] ,
    \top_I.branch[8].l_um_iw[24] ,
    \top_I.branch[8].l_um_iw[23] ,
    \top_I.branch[8].l_um_iw[22] ,
    \top_I.branch[8].l_um_iw[21] ,
    \top_I.branch[8].l_um_iw[20] ,
    \top_I.branch[8].l_um_iw[19] ,
    \top_I.branch[8].l_um_iw[18] ,
    \top_I.branch[8].l_um_iw[17] ,
    \top_I.branch[8].l_um_iw[16] ,
    \top_I.branch[8].l_um_iw[15] ,
    \top_I.branch[8].l_um_iw[14] ,
    \top_I.branch[8].l_um_iw[13] ,
    \top_I.branch[8].l_um_iw[12] ,
    \top_I.branch[8].l_um_iw[11] ,
    \top_I.branch[8].l_um_iw[10] ,
    \top_I.branch[8].l_um_iw[9] ,
    \top_I.branch[8].l_um_iw[8] ,
    \top_I.branch[8].l_um_iw[7] ,
    \top_I.branch[8].l_um_iw[6] ,
    \top_I.branch[8].l_um_iw[5] ,
    \top_I.branch[8].l_um_iw[4] ,
    \top_I.branch[8].l_um_iw[3] ,
    \top_I.branch[8].l_um_iw[2] ,
    \top_I.branch[8].l_um_iw[1] ,
    \top_I.branch[8].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[15] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[14] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[13] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[12] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[11] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[10] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[9] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[8] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[7] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[6] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[5] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[4] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[3] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[2] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].l_um_k_zero[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[8].col_um[0].um_bot_I.uo_out[0] }));
 tt_um_loopback \top_I.branch[9].col_um[0].um_bot_I.block_8_16.tt_um_I  (.clk(\top_I.branch[9].l_um_iw[0] ),
    .ena(\top_I.branch[9].l_um_ena[0] ),
    .rst_n(\top_I.branch[9].l_um_iw[1] ),
    .ui_in({\top_I.branch[9].l_um_iw[9] ,
    \top_I.branch[9].l_um_iw[8] ,
    \top_I.branch[9].l_um_iw[7] ,
    \top_I.branch[9].l_um_iw[6] ,
    \top_I.branch[9].l_um_iw[5] ,
    \top_I.branch[9].l_um_iw[4] ,
    \top_I.branch[9].l_um_iw[3] ,
    \top_I.branch[9].l_um_iw[2] }),
    .uio_in({\top_I.branch[9].l_um_iw[17] ,
    \top_I.branch[9].l_um_iw[16] ,
    \top_I.branch[9].l_um_iw[15] ,
    \top_I.branch[9].l_um_iw[14] ,
    \top_I.branch[9].l_um_iw[13] ,
    \top_I.branch[9].l_um_iw[12] ,
    \top_I.branch[9].l_um_iw[11] ,
    \top_I.branch[9].l_um_iw[10] }),
    .uio_oe({\top_I.branch[9].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[0] }),
    .uio_out({\top_I.branch[9].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[0] }),
    .uo_out({\top_I.branch[9].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[0] }));
 tt_mux \top_I.branch[9].mux_I  (.k_one(\top_I.branch[9].l_k_one ),
    .k_zero(\top_I.branch[9].l_k_zero ),
    .addr({\top_I.branch[9].l_k_zero ,
    \top_I.branch[9].l_k_one ,
    \top_I.branch[9].l_k_zero ,
    \top_I.branch[9].l_k_zero ,
    \top_I.branch[9].l_k_one }),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }),
    .um_ena({\top_I.branch[9].l_um_ena[15] ,
    \top_I.branch[9].l_um_ena[14] ,
    \top_I.branch[9].l_um_ena[13] ,
    \top_I.branch[9].l_um_ena[12] ,
    \top_I.branch[9].l_um_ena[11] ,
    \top_I.branch[9].l_um_ena[10] ,
    \top_I.branch[9].l_um_ena[9] ,
    \top_I.branch[9].l_um_ena[8] ,
    \top_I.branch[9].l_um_ena[7] ,
    \top_I.branch[9].l_um_ena[6] ,
    \top_I.branch[9].l_um_ena[5] ,
    \top_I.branch[9].l_um_ena[4] ,
    \top_I.branch[9].l_um_ena[3] ,
    \top_I.branch[9].l_um_ena[2] ,
    \top_I.branch[9].l_um_ena[1] ,
    \top_I.branch[9].l_um_ena[0] }),
    .um_iw({\top_I.branch[9].l_um_iw[287] ,
    \top_I.branch[9].l_um_iw[286] ,
    \top_I.branch[9].l_um_iw[285] ,
    \top_I.branch[9].l_um_iw[284] ,
    \top_I.branch[9].l_um_iw[283] ,
    \top_I.branch[9].l_um_iw[282] ,
    \top_I.branch[9].l_um_iw[281] ,
    \top_I.branch[9].l_um_iw[280] ,
    \top_I.branch[9].l_um_iw[279] ,
    \top_I.branch[9].l_um_iw[278] ,
    \top_I.branch[9].l_um_iw[277] ,
    \top_I.branch[9].l_um_iw[276] ,
    \top_I.branch[9].l_um_iw[275] ,
    \top_I.branch[9].l_um_iw[274] ,
    \top_I.branch[9].l_um_iw[273] ,
    \top_I.branch[9].l_um_iw[272] ,
    \top_I.branch[9].l_um_iw[271] ,
    \top_I.branch[9].l_um_iw[270] ,
    \top_I.branch[9].l_um_iw[269] ,
    \top_I.branch[9].l_um_iw[268] ,
    \top_I.branch[9].l_um_iw[267] ,
    \top_I.branch[9].l_um_iw[266] ,
    \top_I.branch[9].l_um_iw[265] ,
    \top_I.branch[9].l_um_iw[264] ,
    \top_I.branch[9].l_um_iw[263] ,
    \top_I.branch[9].l_um_iw[262] ,
    \top_I.branch[9].l_um_iw[261] ,
    \top_I.branch[9].l_um_iw[260] ,
    \top_I.branch[9].l_um_iw[259] ,
    \top_I.branch[9].l_um_iw[258] ,
    \top_I.branch[9].l_um_iw[257] ,
    \top_I.branch[9].l_um_iw[256] ,
    \top_I.branch[9].l_um_iw[255] ,
    \top_I.branch[9].l_um_iw[254] ,
    \top_I.branch[9].l_um_iw[253] ,
    \top_I.branch[9].l_um_iw[252] ,
    \top_I.branch[9].l_um_iw[251] ,
    \top_I.branch[9].l_um_iw[250] ,
    \top_I.branch[9].l_um_iw[249] ,
    \top_I.branch[9].l_um_iw[248] ,
    \top_I.branch[9].l_um_iw[247] ,
    \top_I.branch[9].l_um_iw[246] ,
    \top_I.branch[9].l_um_iw[245] ,
    \top_I.branch[9].l_um_iw[244] ,
    \top_I.branch[9].l_um_iw[243] ,
    \top_I.branch[9].l_um_iw[242] ,
    \top_I.branch[9].l_um_iw[241] ,
    \top_I.branch[9].l_um_iw[240] ,
    \top_I.branch[9].l_um_iw[239] ,
    \top_I.branch[9].l_um_iw[238] ,
    \top_I.branch[9].l_um_iw[237] ,
    \top_I.branch[9].l_um_iw[236] ,
    \top_I.branch[9].l_um_iw[235] ,
    \top_I.branch[9].l_um_iw[234] ,
    \top_I.branch[9].l_um_iw[233] ,
    \top_I.branch[9].l_um_iw[232] ,
    \top_I.branch[9].l_um_iw[231] ,
    \top_I.branch[9].l_um_iw[230] ,
    \top_I.branch[9].l_um_iw[229] ,
    \top_I.branch[9].l_um_iw[228] ,
    \top_I.branch[9].l_um_iw[227] ,
    \top_I.branch[9].l_um_iw[226] ,
    \top_I.branch[9].l_um_iw[225] ,
    \top_I.branch[9].l_um_iw[224] ,
    \top_I.branch[9].l_um_iw[223] ,
    \top_I.branch[9].l_um_iw[222] ,
    \top_I.branch[9].l_um_iw[221] ,
    \top_I.branch[9].l_um_iw[220] ,
    \top_I.branch[9].l_um_iw[219] ,
    \top_I.branch[9].l_um_iw[218] ,
    \top_I.branch[9].l_um_iw[217] ,
    \top_I.branch[9].l_um_iw[216] ,
    \top_I.branch[9].l_um_iw[215] ,
    \top_I.branch[9].l_um_iw[214] ,
    \top_I.branch[9].l_um_iw[213] ,
    \top_I.branch[9].l_um_iw[212] ,
    \top_I.branch[9].l_um_iw[211] ,
    \top_I.branch[9].l_um_iw[210] ,
    \top_I.branch[9].l_um_iw[209] ,
    \top_I.branch[9].l_um_iw[208] ,
    \top_I.branch[9].l_um_iw[207] ,
    \top_I.branch[9].l_um_iw[206] ,
    \top_I.branch[9].l_um_iw[205] ,
    \top_I.branch[9].l_um_iw[204] ,
    \top_I.branch[9].l_um_iw[203] ,
    \top_I.branch[9].l_um_iw[202] ,
    \top_I.branch[9].l_um_iw[201] ,
    \top_I.branch[9].l_um_iw[200] ,
    \top_I.branch[9].l_um_iw[199] ,
    \top_I.branch[9].l_um_iw[198] ,
    \top_I.branch[9].l_um_iw[197] ,
    \top_I.branch[9].l_um_iw[196] ,
    \top_I.branch[9].l_um_iw[195] ,
    \top_I.branch[9].l_um_iw[194] ,
    \top_I.branch[9].l_um_iw[193] ,
    \top_I.branch[9].l_um_iw[192] ,
    \top_I.branch[9].l_um_iw[191] ,
    \top_I.branch[9].l_um_iw[190] ,
    \top_I.branch[9].l_um_iw[189] ,
    \top_I.branch[9].l_um_iw[188] ,
    \top_I.branch[9].l_um_iw[187] ,
    \top_I.branch[9].l_um_iw[186] ,
    \top_I.branch[9].l_um_iw[185] ,
    \top_I.branch[9].l_um_iw[184] ,
    \top_I.branch[9].l_um_iw[183] ,
    \top_I.branch[9].l_um_iw[182] ,
    \top_I.branch[9].l_um_iw[181] ,
    \top_I.branch[9].l_um_iw[180] ,
    \top_I.branch[9].l_um_iw[179] ,
    \top_I.branch[9].l_um_iw[178] ,
    \top_I.branch[9].l_um_iw[177] ,
    \top_I.branch[9].l_um_iw[176] ,
    \top_I.branch[9].l_um_iw[175] ,
    \top_I.branch[9].l_um_iw[174] ,
    \top_I.branch[9].l_um_iw[173] ,
    \top_I.branch[9].l_um_iw[172] ,
    \top_I.branch[9].l_um_iw[171] ,
    \top_I.branch[9].l_um_iw[170] ,
    \top_I.branch[9].l_um_iw[169] ,
    \top_I.branch[9].l_um_iw[168] ,
    \top_I.branch[9].l_um_iw[167] ,
    \top_I.branch[9].l_um_iw[166] ,
    \top_I.branch[9].l_um_iw[165] ,
    \top_I.branch[9].l_um_iw[164] ,
    \top_I.branch[9].l_um_iw[163] ,
    \top_I.branch[9].l_um_iw[162] ,
    \top_I.branch[9].l_um_iw[161] ,
    \top_I.branch[9].l_um_iw[160] ,
    \top_I.branch[9].l_um_iw[159] ,
    \top_I.branch[9].l_um_iw[158] ,
    \top_I.branch[9].l_um_iw[157] ,
    \top_I.branch[9].l_um_iw[156] ,
    \top_I.branch[9].l_um_iw[155] ,
    \top_I.branch[9].l_um_iw[154] ,
    \top_I.branch[9].l_um_iw[153] ,
    \top_I.branch[9].l_um_iw[152] ,
    \top_I.branch[9].l_um_iw[151] ,
    \top_I.branch[9].l_um_iw[150] ,
    \top_I.branch[9].l_um_iw[149] ,
    \top_I.branch[9].l_um_iw[148] ,
    \top_I.branch[9].l_um_iw[147] ,
    \top_I.branch[9].l_um_iw[146] ,
    \top_I.branch[9].l_um_iw[145] ,
    \top_I.branch[9].l_um_iw[144] ,
    \top_I.branch[9].l_um_iw[143] ,
    \top_I.branch[9].l_um_iw[142] ,
    \top_I.branch[9].l_um_iw[141] ,
    \top_I.branch[9].l_um_iw[140] ,
    \top_I.branch[9].l_um_iw[139] ,
    \top_I.branch[9].l_um_iw[138] ,
    \top_I.branch[9].l_um_iw[137] ,
    \top_I.branch[9].l_um_iw[136] ,
    \top_I.branch[9].l_um_iw[135] ,
    \top_I.branch[9].l_um_iw[134] ,
    \top_I.branch[9].l_um_iw[133] ,
    \top_I.branch[9].l_um_iw[132] ,
    \top_I.branch[9].l_um_iw[131] ,
    \top_I.branch[9].l_um_iw[130] ,
    \top_I.branch[9].l_um_iw[129] ,
    \top_I.branch[9].l_um_iw[128] ,
    \top_I.branch[9].l_um_iw[127] ,
    \top_I.branch[9].l_um_iw[126] ,
    \top_I.branch[9].l_um_iw[125] ,
    \top_I.branch[9].l_um_iw[124] ,
    \top_I.branch[9].l_um_iw[123] ,
    \top_I.branch[9].l_um_iw[122] ,
    \top_I.branch[9].l_um_iw[121] ,
    \top_I.branch[9].l_um_iw[120] ,
    \top_I.branch[9].l_um_iw[119] ,
    \top_I.branch[9].l_um_iw[118] ,
    \top_I.branch[9].l_um_iw[117] ,
    \top_I.branch[9].l_um_iw[116] ,
    \top_I.branch[9].l_um_iw[115] ,
    \top_I.branch[9].l_um_iw[114] ,
    \top_I.branch[9].l_um_iw[113] ,
    \top_I.branch[9].l_um_iw[112] ,
    \top_I.branch[9].l_um_iw[111] ,
    \top_I.branch[9].l_um_iw[110] ,
    \top_I.branch[9].l_um_iw[109] ,
    \top_I.branch[9].l_um_iw[108] ,
    \top_I.branch[9].l_um_iw[107] ,
    \top_I.branch[9].l_um_iw[106] ,
    \top_I.branch[9].l_um_iw[105] ,
    \top_I.branch[9].l_um_iw[104] ,
    \top_I.branch[9].l_um_iw[103] ,
    \top_I.branch[9].l_um_iw[102] ,
    \top_I.branch[9].l_um_iw[101] ,
    \top_I.branch[9].l_um_iw[100] ,
    \top_I.branch[9].l_um_iw[99] ,
    \top_I.branch[9].l_um_iw[98] ,
    \top_I.branch[9].l_um_iw[97] ,
    \top_I.branch[9].l_um_iw[96] ,
    \top_I.branch[9].l_um_iw[95] ,
    \top_I.branch[9].l_um_iw[94] ,
    \top_I.branch[9].l_um_iw[93] ,
    \top_I.branch[9].l_um_iw[92] ,
    \top_I.branch[9].l_um_iw[91] ,
    \top_I.branch[9].l_um_iw[90] ,
    \top_I.branch[9].l_um_iw[89] ,
    \top_I.branch[9].l_um_iw[88] ,
    \top_I.branch[9].l_um_iw[87] ,
    \top_I.branch[9].l_um_iw[86] ,
    \top_I.branch[9].l_um_iw[85] ,
    \top_I.branch[9].l_um_iw[84] ,
    \top_I.branch[9].l_um_iw[83] ,
    \top_I.branch[9].l_um_iw[82] ,
    \top_I.branch[9].l_um_iw[81] ,
    \top_I.branch[9].l_um_iw[80] ,
    \top_I.branch[9].l_um_iw[79] ,
    \top_I.branch[9].l_um_iw[78] ,
    \top_I.branch[9].l_um_iw[77] ,
    \top_I.branch[9].l_um_iw[76] ,
    \top_I.branch[9].l_um_iw[75] ,
    \top_I.branch[9].l_um_iw[74] ,
    \top_I.branch[9].l_um_iw[73] ,
    \top_I.branch[9].l_um_iw[72] ,
    \top_I.branch[9].l_um_iw[71] ,
    \top_I.branch[9].l_um_iw[70] ,
    \top_I.branch[9].l_um_iw[69] ,
    \top_I.branch[9].l_um_iw[68] ,
    \top_I.branch[9].l_um_iw[67] ,
    \top_I.branch[9].l_um_iw[66] ,
    \top_I.branch[9].l_um_iw[65] ,
    \top_I.branch[9].l_um_iw[64] ,
    \top_I.branch[9].l_um_iw[63] ,
    \top_I.branch[9].l_um_iw[62] ,
    \top_I.branch[9].l_um_iw[61] ,
    \top_I.branch[9].l_um_iw[60] ,
    \top_I.branch[9].l_um_iw[59] ,
    \top_I.branch[9].l_um_iw[58] ,
    \top_I.branch[9].l_um_iw[57] ,
    \top_I.branch[9].l_um_iw[56] ,
    \top_I.branch[9].l_um_iw[55] ,
    \top_I.branch[9].l_um_iw[54] ,
    \top_I.branch[9].l_um_iw[53] ,
    \top_I.branch[9].l_um_iw[52] ,
    \top_I.branch[9].l_um_iw[51] ,
    \top_I.branch[9].l_um_iw[50] ,
    \top_I.branch[9].l_um_iw[49] ,
    \top_I.branch[9].l_um_iw[48] ,
    \top_I.branch[9].l_um_iw[47] ,
    \top_I.branch[9].l_um_iw[46] ,
    \top_I.branch[9].l_um_iw[45] ,
    \top_I.branch[9].l_um_iw[44] ,
    \top_I.branch[9].l_um_iw[43] ,
    \top_I.branch[9].l_um_iw[42] ,
    \top_I.branch[9].l_um_iw[41] ,
    \top_I.branch[9].l_um_iw[40] ,
    \top_I.branch[9].l_um_iw[39] ,
    \top_I.branch[9].l_um_iw[38] ,
    \top_I.branch[9].l_um_iw[37] ,
    \top_I.branch[9].l_um_iw[36] ,
    \top_I.branch[9].l_um_iw[35] ,
    \top_I.branch[9].l_um_iw[34] ,
    \top_I.branch[9].l_um_iw[33] ,
    \top_I.branch[9].l_um_iw[32] ,
    \top_I.branch[9].l_um_iw[31] ,
    \top_I.branch[9].l_um_iw[30] ,
    \top_I.branch[9].l_um_iw[29] ,
    \top_I.branch[9].l_um_iw[28] ,
    \top_I.branch[9].l_um_iw[27] ,
    \top_I.branch[9].l_um_iw[26] ,
    \top_I.branch[9].l_um_iw[25] ,
    \top_I.branch[9].l_um_iw[24] ,
    \top_I.branch[9].l_um_iw[23] ,
    \top_I.branch[9].l_um_iw[22] ,
    \top_I.branch[9].l_um_iw[21] ,
    \top_I.branch[9].l_um_iw[20] ,
    \top_I.branch[9].l_um_iw[19] ,
    \top_I.branch[9].l_um_iw[18] ,
    \top_I.branch[9].l_um_iw[17] ,
    \top_I.branch[9].l_um_iw[16] ,
    \top_I.branch[9].l_um_iw[15] ,
    \top_I.branch[9].l_um_iw[14] ,
    \top_I.branch[9].l_um_iw[13] ,
    \top_I.branch[9].l_um_iw[12] ,
    \top_I.branch[9].l_um_iw[11] ,
    \top_I.branch[9].l_um_iw[10] ,
    \top_I.branch[9].l_um_iw[9] ,
    \top_I.branch[9].l_um_iw[8] ,
    \top_I.branch[9].l_um_iw[7] ,
    \top_I.branch[9].l_um_iw[6] ,
    \top_I.branch[9].l_um_iw[5] ,
    \top_I.branch[9].l_um_iw[4] ,
    \top_I.branch[9].l_um_iw[3] ,
    \top_I.branch[9].l_um_iw[2] ,
    \top_I.branch[9].l_um_iw[1] ,
    \top_I.branch[9].l_um_iw[0] }),
    .um_k_zero({\top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[0] }),
    .um_ow({\top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[15] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[14] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[13] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[12] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[11] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[10] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[9] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[8] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[7] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[6] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[5] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[4] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[3] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[2] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].l_um_k_zero[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_oe[0] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uio_out[0] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[7] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[6] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[5] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[4] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[3] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[2] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[1] ,
    \top_I.branch[9].col_um[0].um_bot_I.uo_out[0] }));
 tt_ctrl \top_I.ctrl_I  (.ctrl_ena(io_in[32]),
    .ctrl_sel_inc(io_in[34]),
    .ctrl_sel_rst_n(io_in[36]),
    .k_one(\top_I.k_one ),
    .k_zero(wbs_ack_o),
    .pad_ui_in({io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6]}),
    .pad_uio_in({io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24]}),
    .pad_uio_oe_n({io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24]}),
    .pad_uio_out({io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24]}),
    .pad_uo_out({io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16]}),
    .spine_iw({\top_I.spine_iw[30] ,
    \top_I.spine_iw[29] ,
    \top_I.spine_iw[28] ,
    \top_I.spine_iw[27] ,
    \top_I.spine_iw[26] ,
    \top_I.spine_iw[25] ,
    \top_I.spine_iw[24] ,
    \top_I.spine_iw[23] ,
    \top_I.spine_iw[22] ,
    \top_I.spine_iw[21] ,
    \top_I.spine_iw[20] ,
    \top_I.spine_iw[19] ,
    \top_I.spine_iw[18] ,
    \top_I.spine_iw[17] ,
    \top_I.spine_iw[16] ,
    \top_I.spine_iw[15] ,
    \top_I.spine_iw[14] ,
    \top_I.spine_iw[13] ,
    \top_I.spine_iw[12] ,
    \top_I.spine_iw[11] ,
    \top_I.spine_iw[10] ,
    \top_I.spine_iw[9] ,
    \top_I.spine_iw[8] ,
    \top_I.spine_iw[7] ,
    \top_I.spine_iw[6] ,
    \top_I.spine_iw[5] ,
    \top_I.spine_iw[4] ,
    \top_I.spine_iw[3] ,
    \top_I.spine_iw[2] ,
    \top_I.spine_iw[1] ,
    \top_I.spine_iw[0] }),
    .spine_ow({\top_I.spine_ow[25] ,
    \top_I.spine_ow[24] ,
    \top_I.spine_ow[23] ,
    \top_I.spine_ow[22] ,
    \top_I.spine_ow[21] ,
    \top_I.spine_ow[20] ,
    \top_I.spine_ow[19] ,
    \top_I.spine_ow[18] ,
    \top_I.spine_ow[17] ,
    \top_I.spine_ow[16] ,
    \top_I.spine_ow[15] ,
    \top_I.spine_ow[14] ,
    \top_I.spine_ow[13] ,
    \top_I.spine_ow[12] ,
    \top_I.spine_ow[11] ,
    \top_I.spine_ow[10] ,
    \top_I.spine_ow[9] ,
    \top_I.spine_ow[8] ,
    \top_I.spine_ow[7] ,
    \top_I.spine_ow[6] ,
    \top_I.spine_ow[5] ,
    \top_I.spine_ow[4] ,
    \top_I.spine_ow[3] ,
    \top_I.spine_ow[2] ,
    \top_I.spine_ow[1] ,
    \top_I.spine_ow[0] }));
 assign io_oeb[0] = \top_I.k_one ;
 assign io_oeb[10] = \top_I.k_one ;
 assign io_oeb[11] = \top_I.k_one ;
 assign io_oeb[12] = \top_I.k_one ;
 assign io_oeb[13] = \top_I.k_one ;
 assign io_oeb[14] = \top_I.k_one ;
 assign io_oeb[15] = \top_I.k_one ;
 assign io_oeb[1] = \top_I.k_one ;
 assign io_oeb[2] = \top_I.k_one ;
 assign io_oeb[32] = \top_I.k_one ;
 assign io_oeb[34] = \top_I.k_one ;
 assign io_oeb[36] = \top_I.k_one ;
 assign io_oeb[3] = \top_I.k_one ;
 assign io_oeb[6] = \top_I.k_one ;
 assign io_oeb[7] = \top_I.k_one ;
 assign io_oeb[8] = \top_I.k_one ;
 assign io_oeb[9] = \top_I.k_one ;
 assign io_out[0] = \top_I.k_one ;
 assign io_out[10] = \top_I.k_one ;
 assign io_out[11] = \top_I.k_one ;
 assign io_out[12] = \top_I.k_one ;
 assign io_out[13] = \top_I.k_one ;
 assign io_out[14] = \top_I.k_one ;
 assign io_out[15] = \top_I.k_one ;
 assign io_out[1] = \top_I.k_one ;
 assign io_out[2] = \top_I.k_one ;
 assign io_out[3] = \top_I.k_one ;
 assign io_out[6] = \top_I.k_one ;
 assign io_out[7] = \top_I.k_one ;
 assign io_out[8] = \top_I.k_one ;
 assign io_out[9] = \top_I.k_one ;
 assign io_out[5] = user_clock2;
 assign io_oeb[16] = wbs_ack_o;
 assign io_oeb[17] = wbs_ack_o;
 assign io_oeb[18] = wbs_ack_o;
 assign io_oeb[19] = wbs_ack_o;
 assign io_oeb[20] = wbs_ack_o;
 assign io_oeb[21] = wbs_ack_o;
 assign io_oeb[22] = wbs_ack_o;
 assign io_oeb[23] = wbs_ack_o;
 assign io_oeb[33] = wbs_ack_o;
 assign io_oeb[35] = wbs_ack_o;
 assign io_oeb[37] = wbs_ack_o;
 assign io_oeb[4] = wbs_ack_o;
 assign io_oeb[5] = wbs_ack_o;
 assign io_out[32] = wbs_ack_o;
 assign io_out[33] = wbs_ack_o;
 assign io_out[34] = wbs_ack_o;
 assign io_out[35] = wbs_ack_o;
 assign io_out[36] = wbs_ack_o;
 assign io_out[37] = wbs_ack_o;
 assign io_out[4] = wbs_ack_o;
 assign la_data_out[0] = wbs_ack_o;
 assign la_data_out[100] = wbs_ack_o;
 assign la_data_out[101] = wbs_ack_o;
 assign la_data_out[102] = wbs_ack_o;
 assign la_data_out[103] = wbs_ack_o;
 assign la_data_out[104] = wbs_ack_o;
 assign la_data_out[105] = wbs_ack_o;
 assign la_data_out[106] = wbs_ack_o;
 assign la_data_out[107] = wbs_ack_o;
 assign la_data_out[108] = wbs_ack_o;
 assign la_data_out[109] = wbs_ack_o;
 assign la_data_out[10] = wbs_ack_o;
 assign la_data_out[110] = wbs_ack_o;
 assign la_data_out[111] = wbs_ack_o;
 assign la_data_out[112] = wbs_ack_o;
 assign la_data_out[113] = wbs_ack_o;
 assign la_data_out[114] = wbs_ack_o;
 assign la_data_out[115] = wbs_ack_o;
 assign la_data_out[116] = wbs_ack_o;
 assign la_data_out[117] = wbs_ack_o;
 assign la_data_out[118] = wbs_ack_o;
 assign la_data_out[119] = wbs_ack_o;
 assign la_data_out[11] = wbs_ack_o;
 assign la_data_out[120] = wbs_ack_o;
 assign la_data_out[121] = wbs_ack_o;
 assign la_data_out[122] = wbs_ack_o;
 assign la_data_out[123] = wbs_ack_o;
 assign la_data_out[124] = wbs_ack_o;
 assign la_data_out[125] = wbs_ack_o;
 assign la_data_out[126] = wbs_ack_o;
 assign la_data_out[127] = wbs_ack_o;
 assign la_data_out[12] = wbs_ack_o;
 assign la_data_out[13] = wbs_ack_o;
 assign la_data_out[14] = wbs_ack_o;
 assign la_data_out[15] = wbs_ack_o;
 assign la_data_out[16] = wbs_ack_o;
 assign la_data_out[17] = wbs_ack_o;
 assign la_data_out[18] = wbs_ack_o;
 assign la_data_out[19] = wbs_ack_o;
 assign la_data_out[1] = wbs_ack_o;
 assign la_data_out[20] = wbs_ack_o;
 assign la_data_out[21] = wbs_ack_o;
 assign la_data_out[22] = wbs_ack_o;
 assign la_data_out[23] = wbs_ack_o;
 assign la_data_out[24] = wbs_ack_o;
 assign la_data_out[25] = wbs_ack_o;
 assign la_data_out[26] = wbs_ack_o;
 assign la_data_out[27] = wbs_ack_o;
 assign la_data_out[28] = wbs_ack_o;
 assign la_data_out[29] = wbs_ack_o;
 assign la_data_out[2] = wbs_ack_o;
 assign la_data_out[30] = wbs_ack_o;
 assign la_data_out[31] = wbs_ack_o;
 assign la_data_out[32] = wbs_ack_o;
 assign la_data_out[33] = wbs_ack_o;
 assign la_data_out[34] = wbs_ack_o;
 assign la_data_out[35] = wbs_ack_o;
 assign la_data_out[36] = wbs_ack_o;
 assign la_data_out[37] = wbs_ack_o;
 assign la_data_out[38] = wbs_ack_o;
 assign la_data_out[39] = wbs_ack_o;
 assign la_data_out[3] = wbs_ack_o;
 assign la_data_out[40] = wbs_ack_o;
 assign la_data_out[41] = wbs_ack_o;
 assign la_data_out[42] = wbs_ack_o;
 assign la_data_out[43] = wbs_ack_o;
 assign la_data_out[44] = wbs_ack_o;
 assign la_data_out[45] = wbs_ack_o;
 assign la_data_out[46] = wbs_ack_o;
 assign la_data_out[47] = wbs_ack_o;
 assign la_data_out[48] = wbs_ack_o;
 assign la_data_out[49] = wbs_ack_o;
 assign la_data_out[4] = wbs_ack_o;
 assign la_data_out[50] = wbs_ack_o;
 assign la_data_out[51] = wbs_ack_o;
 assign la_data_out[52] = wbs_ack_o;
 assign la_data_out[53] = wbs_ack_o;
 assign la_data_out[54] = wbs_ack_o;
 assign la_data_out[55] = wbs_ack_o;
 assign la_data_out[56] = wbs_ack_o;
 assign la_data_out[57] = wbs_ack_o;
 assign la_data_out[58] = wbs_ack_o;
 assign la_data_out[59] = wbs_ack_o;
 assign la_data_out[5] = wbs_ack_o;
 assign la_data_out[60] = wbs_ack_o;
 assign la_data_out[61] = wbs_ack_o;
 assign la_data_out[62] = wbs_ack_o;
 assign la_data_out[63] = wbs_ack_o;
 assign la_data_out[64] = wbs_ack_o;
 assign la_data_out[65] = wbs_ack_o;
 assign la_data_out[66] = wbs_ack_o;
 assign la_data_out[67] = wbs_ack_o;
 assign la_data_out[68] = wbs_ack_o;
 assign la_data_out[69] = wbs_ack_o;
 assign la_data_out[6] = wbs_ack_o;
 assign la_data_out[70] = wbs_ack_o;
 assign la_data_out[71] = wbs_ack_o;
 assign la_data_out[72] = wbs_ack_o;
 assign la_data_out[73] = wbs_ack_o;
 assign la_data_out[74] = wbs_ack_o;
 assign la_data_out[75] = wbs_ack_o;
 assign la_data_out[76] = wbs_ack_o;
 assign la_data_out[77] = wbs_ack_o;
 assign la_data_out[78] = wbs_ack_o;
 assign la_data_out[79] = wbs_ack_o;
 assign la_data_out[7] = wbs_ack_o;
 assign la_data_out[80] = wbs_ack_o;
 assign la_data_out[81] = wbs_ack_o;
 assign la_data_out[82] = wbs_ack_o;
 assign la_data_out[83] = wbs_ack_o;
 assign la_data_out[84] = wbs_ack_o;
 assign la_data_out[85] = wbs_ack_o;
 assign la_data_out[86] = wbs_ack_o;
 assign la_data_out[87] = wbs_ack_o;
 assign la_data_out[88] = wbs_ack_o;
 assign la_data_out[89] = wbs_ack_o;
 assign la_data_out[8] = wbs_ack_o;
 assign la_data_out[90] = wbs_ack_o;
 assign la_data_out[91] = wbs_ack_o;
 assign la_data_out[92] = wbs_ack_o;
 assign la_data_out[93] = wbs_ack_o;
 assign la_data_out[94] = wbs_ack_o;
 assign la_data_out[95] = wbs_ack_o;
 assign la_data_out[96] = wbs_ack_o;
 assign la_data_out[97] = wbs_ack_o;
 assign la_data_out[98] = wbs_ack_o;
 assign la_data_out[99] = wbs_ack_o;
 assign la_data_out[9] = wbs_ack_o;
 assign user_irq[0] = wbs_ack_o;
 assign user_irq[1] = wbs_ack_o;
 assign user_irq[2] = wbs_ack_o;
 assign wbs_dat_o[0] = wbs_ack_o;
 assign wbs_dat_o[10] = wbs_ack_o;
 assign wbs_dat_o[11] = wbs_ack_o;
 assign wbs_dat_o[12] = wbs_ack_o;
 assign wbs_dat_o[13] = wbs_ack_o;
 assign wbs_dat_o[14] = wbs_ack_o;
 assign wbs_dat_o[15] = wbs_ack_o;
 assign wbs_dat_o[16] = wbs_ack_o;
 assign wbs_dat_o[17] = wbs_ack_o;
 assign wbs_dat_o[18] = wbs_ack_o;
 assign wbs_dat_o[19] = wbs_ack_o;
 assign wbs_dat_o[1] = wbs_ack_o;
 assign wbs_dat_o[20] = wbs_ack_o;
 assign wbs_dat_o[21] = wbs_ack_o;
 assign wbs_dat_o[22] = wbs_ack_o;
 assign wbs_dat_o[23] = wbs_ack_o;
 assign wbs_dat_o[24] = wbs_ack_o;
 assign wbs_dat_o[25] = wbs_ack_o;
 assign wbs_dat_o[26] = wbs_ack_o;
 assign wbs_dat_o[27] = wbs_ack_o;
 assign wbs_dat_o[28] = wbs_ack_o;
 assign wbs_dat_o[29] = wbs_ack_o;
 assign wbs_dat_o[2] = wbs_ack_o;
 assign wbs_dat_o[30] = wbs_ack_o;
 assign wbs_dat_o[31] = wbs_ack_o;
 assign wbs_dat_o[3] = wbs_ack_o;
 assign wbs_dat_o[4] = wbs_ack_o;
 assign wbs_dat_o[5] = wbs_ack_o;
 assign wbs_dat_o[6] = wbs_ack_o;
 assign wbs_dat_o[7] = wbs_ack_o;
 assign wbs_dat_o[8] = wbs_ack_o;
 assign wbs_dat_o[9] = wbs_ack_o;
endmodule
