VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_as1802
  CLASS BLOCK ;
  FOREIGN tt_um_as1802 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1362.520 BY 220.320 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 219.150 158.850 220.320 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 219.320 162.530 220.320 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 218.100 155.170 220.320 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 216.740 151.490 220.320 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 215.380 147.810 220.320 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 216.740 144.130 220.320 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 215.380 140.450 220.320 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 215.380 136.770 220.320 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 216.740 133.090 220.320 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 216.740 129.410 220.320 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 219.320 125.730 220.320 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 214.020 122.050 220.320 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 214.020 118.370 220.320 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 218.100 114.690 220.320 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 218.780 111.010 220.320 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 218.780 107.330 220.320 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 211.300 103.650 220.320 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 216.060 99.970 220.320 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 218.780 96.290 220.320 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 218.100 33.730 220.320 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 218.780 30.050 220.320 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 218.780 26.370 220.320 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 218.100 22.690 220.320 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 218.100 19.010 220.320 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 218.780 15.330 220.320 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 218.780 11.650 220.320 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 218.780 7.970 220.320 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 193.620 63.170 220.320 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 199.740 59.490 220.320 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 193.620 55.810 220.320 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 194.980 52.130 220.320 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 195.660 48.450 220.320 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 193.620 44.770 220.320 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 193.620 41.090 220.320 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 194.300 37.410 220.320 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 193.620 92.610 220.320 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 214.700 88.930 220.320 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 218.780 85.250 220.320 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 218.780 81.570 220.320 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 193.620 77.890 220.320 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 218.780 74.210 220.320 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 218.780 70.530 220.320 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 218.780 66.850 220.320 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 5.200 329.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 5.200 483.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 5.200 637.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 5.200 790.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 5.200 944.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 5.200 1097.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 5.200 1251.440 215.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 5.200 253.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 5.200 406.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 5.200 560.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 5.200 713.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 5.200 867.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 5.200 1021.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 5.200 1174.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 5.200 1328.240 215.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 213.465 1357.190 215.070 ;
        RECT 5.330 208.025 1357.190 210.855 ;
        RECT 5.330 202.585 1357.190 205.415 ;
        RECT 5.330 197.145 1357.190 199.975 ;
        RECT 5.330 191.705 1357.190 194.535 ;
        RECT 5.330 186.265 1357.190 189.095 ;
        RECT 5.330 180.825 1357.190 183.655 ;
        RECT 5.330 175.385 1357.190 178.215 ;
        RECT 5.330 169.945 1357.190 172.775 ;
        RECT 5.330 164.505 1357.190 167.335 ;
        RECT 5.330 159.065 1357.190 161.895 ;
        RECT 5.330 153.625 1357.190 156.455 ;
        RECT 5.330 148.185 1357.190 151.015 ;
        RECT 5.330 142.745 1357.190 145.575 ;
        RECT 5.330 137.305 1357.190 140.135 ;
        RECT 5.330 131.865 1357.190 134.695 ;
        RECT 5.330 126.425 1357.190 129.255 ;
        RECT 5.330 120.985 1357.190 123.815 ;
        RECT 5.330 115.545 1357.190 118.375 ;
        RECT 5.330 110.105 1357.190 112.935 ;
        RECT 5.330 104.665 1357.190 107.495 ;
        RECT 5.330 99.225 1357.190 102.055 ;
        RECT 5.330 93.785 1357.190 96.615 ;
        RECT 5.330 88.345 1357.190 91.175 ;
        RECT 5.330 82.905 1357.190 85.735 ;
        RECT 5.330 77.465 1357.190 80.295 ;
        RECT 5.330 72.025 1357.190 74.855 ;
        RECT 5.330 66.585 1357.190 69.415 ;
        RECT 5.330 61.145 1357.190 63.975 ;
        RECT 5.330 55.705 1357.190 58.535 ;
        RECT 5.330 50.265 1357.190 53.095 ;
        RECT 5.330 44.825 1357.190 47.655 ;
        RECT 5.330 39.385 1357.190 42.215 ;
        RECT 5.330 33.945 1357.190 36.775 ;
        RECT 5.330 28.505 1357.190 31.335 ;
        RECT 5.330 23.065 1357.190 25.895 ;
        RECT 5.330 17.625 1357.190 20.455 ;
        RECT 5.330 12.185 1357.190 15.015 ;
        RECT 5.330 6.745 1357.190 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 1357.000 214.965 ;
      LAYER met1 ;
        RECT 5.520 0.040 1357.000 220.280 ;
      LAYER met2 ;
        RECT 10.670 0.010 1344.940 220.310 ;
      LAYER met3 ;
        RECT 7.630 0.175 1340.375 220.145 ;
      LAYER met4 ;
        RECT 8.370 218.380 10.950 220.145 ;
        RECT 12.050 218.380 14.630 220.145 ;
        RECT 15.730 218.380 18.310 220.145 ;
        RECT 7.655 217.700 18.310 218.380 ;
        RECT 19.410 217.700 21.990 220.145 ;
        RECT 23.090 218.380 25.670 220.145 ;
        RECT 26.770 218.380 29.350 220.145 ;
        RECT 30.450 218.380 33.030 220.145 ;
        RECT 23.090 217.700 33.030 218.380 ;
        RECT 34.130 217.700 36.710 220.145 ;
        RECT 7.655 215.520 36.710 217.700 ;
        RECT 7.655 4.800 20.640 215.520 ;
        RECT 23.040 193.900 36.710 215.520 ;
        RECT 37.810 193.900 40.390 220.145 ;
        RECT 23.040 193.220 40.390 193.900 ;
        RECT 41.490 193.220 44.070 220.145 ;
        RECT 45.170 195.260 47.750 220.145 ;
        RECT 48.850 195.260 51.430 220.145 ;
        RECT 45.170 194.580 51.430 195.260 ;
        RECT 52.530 194.580 55.110 220.145 ;
        RECT 45.170 193.220 55.110 194.580 ;
        RECT 56.210 199.340 58.790 220.145 ;
        RECT 59.890 199.340 62.470 220.145 ;
        RECT 56.210 193.220 62.470 199.340 ;
        RECT 63.570 218.380 66.150 220.145 ;
        RECT 67.250 218.380 69.830 220.145 ;
        RECT 70.930 218.380 73.510 220.145 ;
        RECT 74.610 218.380 77.190 220.145 ;
        RECT 63.570 193.220 77.190 218.380 ;
        RECT 78.290 218.380 80.870 220.145 ;
        RECT 81.970 218.380 84.550 220.145 ;
        RECT 85.650 218.380 88.230 220.145 ;
        RECT 78.290 214.300 88.230 218.380 ;
        RECT 89.330 214.300 91.910 220.145 ;
        RECT 78.290 193.220 91.910 214.300 ;
        RECT 93.010 218.380 95.590 220.145 ;
        RECT 96.690 218.380 99.270 220.145 ;
        RECT 93.010 215.660 99.270 218.380 ;
        RECT 100.370 215.660 102.950 220.145 ;
        RECT 93.010 215.520 102.950 215.660 ;
        RECT 93.010 193.220 97.440 215.520 ;
        RECT 23.040 4.800 97.440 193.220 ;
        RECT 99.840 210.900 102.950 215.520 ;
        RECT 104.050 218.380 106.630 220.145 ;
        RECT 107.730 218.380 110.310 220.145 ;
        RECT 111.410 218.380 113.990 220.145 ;
        RECT 104.050 217.700 113.990 218.380 ;
        RECT 115.090 217.700 117.670 220.145 ;
        RECT 104.050 213.620 117.670 217.700 ;
        RECT 118.770 213.620 121.350 220.145 ;
        RECT 122.450 218.920 125.030 220.145 ;
        RECT 126.130 218.920 128.710 220.145 ;
        RECT 122.450 216.340 128.710 218.920 ;
        RECT 129.810 216.340 132.390 220.145 ;
        RECT 133.490 216.340 136.070 220.145 ;
        RECT 122.450 214.980 136.070 216.340 ;
        RECT 137.170 214.980 139.750 220.145 ;
        RECT 140.850 216.340 143.430 220.145 ;
        RECT 144.530 216.340 147.110 220.145 ;
        RECT 140.850 214.980 147.110 216.340 ;
        RECT 148.210 216.340 150.790 220.145 ;
        RECT 151.890 217.700 154.470 220.145 ;
        RECT 155.570 218.750 158.150 220.145 ;
        RECT 159.250 218.920 161.830 220.145 ;
        RECT 162.930 218.920 1095.425 220.145 ;
        RECT 159.250 218.750 1095.425 218.920 ;
        RECT 155.570 217.700 1095.425 218.750 ;
        RECT 151.890 216.340 1095.425 217.700 ;
        RECT 148.210 215.520 1095.425 216.340 ;
        RECT 148.210 214.980 174.240 215.520 ;
        RECT 122.450 213.620 174.240 214.980 ;
        RECT 104.050 210.900 174.240 213.620 ;
        RECT 99.840 4.800 174.240 210.900 ;
        RECT 176.640 4.800 251.040 215.520 ;
        RECT 253.440 4.800 327.840 215.520 ;
        RECT 330.240 4.800 404.640 215.520 ;
        RECT 407.040 4.800 481.440 215.520 ;
        RECT 483.840 4.800 558.240 215.520 ;
        RECT 560.640 4.800 635.040 215.520 ;
        RECT 637.440 4.800 711.840 215.520 ;
        RECT 714.240 4.800 788.640 215.520 ;
        RECT 791.040 4.800 865.440 215.520 ;
        RECT 867.840 4.800 942.240 215.520 ;
        RECT 944.640 4.800 1019.040 215.520 ;
        RECT 1021.440 4.800 1095.425 215.520 ;
        RECT 7.655 1.535 1095.425 4.800 ;
  END
END tt_um_as1802
END LIBRARY

