VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_mux
  CLASS BLOCK ;
  FOREIGN tt_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 1358.840 BY 54.400 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.480 2.480 711.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.080 2.480 864.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1016.680 2.480 1018.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1170.280 2.480 1171.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.880 2.480 1325.480 51.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.680 2.480 634.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.280 2.480 787.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 939.880 2.480 941.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1093.480 2.480 1095.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1247.080 2.480 1248.680 51.920 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 47.790 1358.840 48.090 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.561000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 47.110 1358.840 47.410 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.493500 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 46.430 1358.840 46.730 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.561000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 45.750 1358.840 46.050 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 45.070 1358.840 45.370 ;
    END
  END addr[4]
  PIN k_one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 44.390 1358.840 44.690 ;
    END
  END k_one
  PIN k_zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 43.710 1358.840 44.010 ;
    END
  END k_zero
  PIN spine_iw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 43.030 1358.840 43.330 ;
    END
  END spine_iw[0]
  PIN spine_iw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.561000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 36.230 1358.840 36.530 ;
    END
  END spine_iw[10]
  PIN spine_iw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.493500 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 35.550 1358.840 35.850 ;
    END
  END spine_iw[11]
  PIN spine_iw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 34.870 1358.840 35.170 ;
    END
  END spine_iw[12]
  PIN spine_iw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 34.190 1358.840 34.490 ;
    END
  END spine_iw[13]
  PIN spine_iw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 33.510 1358.840 33.810 ;
    END
  END spine_iw[14]
  PIN spine_iw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 32.830 1358.840 33.130 ;
    END
  END spine_iw[15]
  PIN spine_iw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 32.150 1358.840 32.450 ;
    END
  END spine_iw[16]
  PIN spine_iw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 31.470 1358.840 31.770 ;
    END
  END spine_iw[17]
  PIN spine_iw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 30.790 1358.840 31.090 ;
    END
  END spine_iw[18]
  PIN spine_iw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 30.110 1358.840 30.410 ;
    END
  END spine_iw[19]
  PIN spine_iw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 42.350 1358.840 42.650 ;
    END
  END spine_iw[1]
  PIN spine_iw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 29.430 1358.840 29.730 ;
    END
  END spine_iw[20]
  PIN spine_iw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 28.750 1358.840 29.050 ;
    END
  END spine_iw[21]
  PIN spine_iw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 28.070 1358.840 28.370 ;
    END
  END spine_iw[22]
  PIN spine_iw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 27.390 1358.840 27.690 ;
    END
  END spine_iw[23]
  PIN spine_iw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 26.710 1358.840 27.010 ;
    END
  END spine_iw[24]
  PIN spine_iw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 26.030 1358.840 26.330 ;
    END
  END spine_iw[25]
  PIN spine_iw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 25.350 1358.840 25.650 ;
    END
  END spine_iw[26]
  PIN spine_iw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 24.670 1358.840 24.970 ;
    END
  END spine_iw[27]
  PIN spine_iw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 23.990 1358.840 24.290 ;
    END
  END spine_iw[28]
  PIN spine_iw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 23.310 1358.840 23.610 ;
    END
  END spine_iw[29]
  PIN spine_iw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 41.670 1358.840 41.970 ;
    END
  END spine_iw[2]
  PIN spine_iw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 22.630 1358.840 22.930 ;
    END
  END spine_iw[30]
  PIN spine_iw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 40.990 1358.840 41.290 ;
    END
  END spine_iw[3]
  PIN spine_iw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 40.310 1358.840 40.610 ;
    END
  END spine_iw[4]
  PIN spine_iw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 39.630 1358.840 39.930 ;
    END
  END spine_iw[5]
  PIN spine_iw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 38.950 1358.840 39.250 ;
    END
  END spine_iw[6]
  PIN spine_iw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 38.270 1358.840 38.570 ;
    END
  END spine_iw[7]
  PIN spine_iw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.561000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 37.590 1358.840 37.890 ;
    END
  END spine_iw[8]
  PIN spine_iw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 36.910 1358.840 37.210 ;
    END
  END spine_iw[9]
  PIN spine_ow[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 21.950 1358.840 22.250 ;
    END
  END spine_ow[0]
  PIN spine_ow[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 15.150 1358.840 15.450 ;
    END
  END spine_ow[10]
  PIN spine_ow[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 14.470 1358.840 14.770 ;
    END
  END spine_ow[11]
  PIN spine_ow[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 13.790 1358.840 14.090 ;
    END
  END spine_ow[12]
  PIN spine_ow[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 13.110 1358.840 13.410 ;
    END
  END spine_ow[13]
  PIN spine_ow[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 12.430 1358.840 12.730 ;
    END
  END spine_ow[14]
  PIN spine_ow[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 11.750 1358.840 12.050 ;
    END
  END spine_ow[15]
  PIN spine_ow[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 11.070 1358.840 11.370 ;
    END
  END spine_ow[16]
  PIN spine_ow[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 10.390 1358.840 10.690 ;
    END
  END spine_ow[17]
  PIN spine_ow[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 9.710 1358.840 10.010 ;
    END
  END spine_ow[18]
  PIN spine_ow[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 9.030 1358.840 9.330 ;
    END
  END spine_ow[19]
  PIN spine_ow[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 21.270 1358.840 21.570 ;
    END
  END spine_ow[1]
  PIN spine_ow[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 8.350 1358.840 8.650 ;
    END
  END spine_ow[20]
  PIN spine_ow[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 7.670 1358.840 7.970 ;
    END
  END spine_ow[21]
  PIN spine_ow[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 6.990 1358.840 7.290 ;
    END
  END spine_ow[22]
  PIN spine_ow[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 6.310 1358.840 6.610 ;
    END
  END spine_ow[23]
  PIN spine_ow[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 5.630 1358.840 5.930 ;
    END
  END spine_ow[24]
  PIN spine_ow[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.840 4.950 1358.840 5.250 ;
    END
  END spine_ow[25]
  PIN spine_ow[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 20.590 1358.840 20.890 ;
    END
  END spine_ow[2]
  PIN spine_ow[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 19.910 1358.840 20.210 ;
    END
  END spine_ow[3]
  PIN spine_ow[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 19.230 1358.840 19.530 ;
    END
  END spine_ow[4]
  PIN spine_ow[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 18.550 1358.840 18.850 ;
    END
  END spine_ow[5]
  PIN spine_ow[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 17.870 1358.840 18.170 ;
    END
  END spine_ow[6]
  PIN spine_ow[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 17.190 1358.840 17.490 ;
    END
  END spine_ow[7]
  PIN spine_ow[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 16.510 1358.840 16.810 ;
    END
  END spine_ow[8]
  PIN spine_ow[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1357.840 15.830 1358.840 16.130 ;
    END
  END spine_ow[9]
  PIN um_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 162.230 0.000 162.530 1.000 ;
    END
  END um_ena[0]
  PIN um_ena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1013.230 0.000 1013.530 1.000 ;
    END
  END um_ena[10]
  PIN um_ena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1013.230 53.400 1013.530 54.400 ;
    END
  END um_ena[11]
  PIN um_ena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1183.430 0.000 1183.730 1.000 ;
    END
  END um_ena[12]
  PIN um_ena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1183.430 53.400 1183.730 54.400 ;
    END
  END um_ena[13]
  PIN um_ena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1353.630 0.000 1353.930 1.000 ;
    END
  END um_ena[14]
  PIN um_ena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1353.630 53.400 1353.930 54.400 ;
    END
  END um_ena[15]
  PIN um_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 162.230 53.400 162.530 54.400 ;
    END
  END um_ena[1]
  PIN um_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 332.430 0.000 332.730 1.000 ;
    END
  END um_ena[2]
  PIN um_ena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 332.430 53.400 332.730 54.400 ;
    END
  END um_ena[3]
  PIN um_ena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 502.630 0.000 502.930 1.000 ;
    END
  END um_ena[4]
  PIN um_ena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 502.630 53.400 502.930 54.400 ;
    END
  END um_ena[5]
  PIN um_ena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 672.830 0.000 673.130 1.000 ;
    END
  END um_ena[6]
  PIN um_ena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 672.830 53.400 673.130 54.400 ;
    END
  END um_ena[7]
  PIN um_ena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 843.030 0.000 843.330 1.000 ;
    END
  END um_ena[8]
  PIN um_ena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 843.030 53.400 843.330 54.400 ;
    END
  END um_ena[9]
  PIN um_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 158.550 0.000 158.850 1.000 ;
    END
  END um_iw[0]
  PIN um_iw[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 462.150 53.400 462.450 54.400 ;
    END
  END um_iw[100]
  PIN um_iw[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 458.470 53.400 458.770 54.400 ;
    END
  END um_iw[101]
  PIN um_iw[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 454.790 53.400 455.090 54.400 ;
    END
  END um_iw[102]
  PIN um_iw[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 451.110 53.400 451.410 54.400 ;
    END
  END um_iw[103]
  PIN um_iw[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 447.430 53.400 447.730 54.400 ;
    END
  END um_iw[104]
  PIN um_iw[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 443.750 53.400 444.050 54.400 ;
    END
  END um_iw[105]
  PIN um_iw[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 440.070 53.400 440.370 54.400 ;
    END
  END um_iw[106]
  PIN um_iw[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 436.390 53.400 436.690 54.400 ;
    END
  END um_iw[107]
  PIN um_iw[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 669.150 0.000 669.450 1.000 ;
    END
  END um_iw[108]
  PIN um_iw[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 665.470 0.000 665.770 1.000 ;
    END
  END um_iw[109]
  PIN um_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 0.000 122.050 1.000 ;
    END
  END um_iw[10]
  PIN um_iw[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 661.790 0.000 662.090 1.000 ;
    END
  END um_iw[110]
  PIN um_iw[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 658.110 0.000 658.410 1.000 ;
    END
  END um_iw[111]
  PIN um_iw[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 654.430 0.000 654.730 1.000 ;
    END
  END um_iw[112]
  PIN um_iw[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 650.750 0.000 651.050 1.000 ;
    END
  END um_iw[113]
  PIN um_iw[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 647.070 0.000 647.370 1.000 ;
    END
  END um_iw[114]
  PIN um_iw[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 643.390 0.000 643.690 1.000 ;
    END
  END um_iw[115]
  PIN um_iw[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 639.710 0.000 640.010 1.000 ;
    END
  END um_iw[116]
  PIN um_iw[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 636.030 0.000 636.330 1.000 ;
    END
  END um_iw[117]
  PIN um_iw[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 632.350 0.000 632.650 1.000 ;
    END
  END um_iw[118]
  PIN um_iw[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 628.670 0.000 628.970 1.000 ;
    END
  END um_iw[119]
  PIN um_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 0.000 118.370 1.000 ;
    END
  END um_iw[11]
  PIN um_iw[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 624.990 0.000 625.290 1.000 ;
    END
  END um_iw[120]
  PIN um_iw[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 621.310 0.000 621.610 1.000 ;
    END
  END um_iw[121]
  PIN um_iw[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 617.630 0.000 617.930 1.000 ;
    END
  END um_iw[122]
  PIN um_iw[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 613.950 0.000 614.250 1.000 ;
    END
  END um_iw[123]
  PIN um_iw[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 610.270 0.000 610.570 1.000 ;
    END
  END um_iw[124]
  PIN um_iw[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 606.590 0.000 606.890 1.000 ;
    END
  END um_iw[125]
  PIN um_iw[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 669.150 53.400 669.450 54.400 ;
    END
  END um_iw[126]
  PIN um_iw[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 665.470 53.400 665.770 54.400 ;
    END
  END um_iw[127]
  PIN um_iw[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 661.790 53.400 662.090 54.400 ;
    END
  END um_iw[128]
  PIN um_iw[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 658.110 53.400 658.410 54.400 ;
    END
  END um_iw[129]
  PIN um_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 0.000 114.690 1.000 ;
    END
  END um_iw[12]
  PIN um_iw[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 654.430 53.400 654.730 54.400 ;
    END
  END um_iw[130]
  PIN um_iw[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 650.750 53.400 651.050 54.400 ;
    END
  END um_iw[131]
  PIN um_iw[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 647.070 53.400 647.370 54.400 ;
    END
  END um_iw[132]
  PIN um_iw[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 643.390 53.400 643.690 54.400 ;
    END
  END um_iw[133]
  PIN um_iw[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 639.710 53.400 640.010 54.400 ;
    END
  END um_iw[134]
  PIN um_iw[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 636.030 53.400 636.330 54.400 ;
    END
  END um_iw[135]
  PIN um_iw[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 632.350 53.400 632.650 54.400 ;
    END
  END um_iw[136]
  PIN um_iw[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 628.670 53.400 628.970 54.400 ;
    END
  END um_iw[137]
  PIN um_iw[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 624.990 53.400 625.290 54.400 ;
    END
  END um_iw[138]
  PIN um_iw[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 621.310 53.400 621.610 54.400 ;
    END
  END um_iw[139]
  PIN um_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 0.000 111.010 1.000 ;
    END
  END um_iw[13]
  PIN um_iw[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 617.630 53.400 617.930 54.400 ;
    END
  END um_iw[140]
  PIN um_iw[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 613.950 53.400 614.250 54.400 ;
    END
  END um_iw[141]
  PIN um_iw[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 610.270 53.400 610.570 54.400 ;
    END
  END um_iw[142]
  PIN um_iw[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 606.590 53.400 606.890 54.400 ;
    END
  END um_iw[143]
  PIN um_iw[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 839.350 0.000 839.650 1.000 ;
    END
  END um_iw[144]
  PIN um_iw[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 835.670 0.000 835.970 1.000 ;
    END
  END um_iw[145]
  PIN um_iw[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 831.990 0.000 832.290 1.000 ;
    END
  END um_iw[146]
  PIN um_iw[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 828.310 0.000 828.610 1.000 ;
    END
  END um_iw[147]
  PIN um_iw[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 824.630 0.000 824.930 1.000 ;
    END
  END um_iw[148]
  PIN um_iw[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 820.950 0.000 821.250 1.000 ;
    END
  END um_iw[149]
  PIN um_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 0.000 107.330 1.000 ;
    END
  END um_iw[14]
  PIN um_iw[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 817.270 0.000 817.570 1.000 ;
    END
  END um_iw[150]
  PIN um_iw[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 813.590 0.000 813.890 1.000 ;
    END
  END um_iw[151]
  PIN um_iw[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 809.910 0.000 810.210 1.000 ;
    END
  END um_iw[152]
  PIN um_iw[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 806.230 0.000 806.530 1.000 ;
    END
  END um_iw[153]
  PIN um_iw[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 802.550 0.000 802.850 1.000 ;
    END
  END um_iw[154]
  PIN um_iw[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 798.870 0.000 799.170 1.000 ;
    END
  END um_iw[155]
  PIN um_iw[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 795.190 0.000 795.490 1.000 ;
    END
  END um_iw[156]
  PIN um_iw[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 791.510 0.000 791.810 1.000 ;
    END
  END um_iw[157]
  PIN um_iw[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 787.830 0.000 788.130 1.000 ;
    END
  END um_iw[158]
  PIN um_iw[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 784.150 0.000 784.450 1.000 ;
    END
  END um_iw[159]
  PIN um_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 103.350 0.000 103.650 1.000 ;
    END
  END um_iw[15]
  PIN um_iw[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 780.470 0.000 780.770 1.000 ;
    END
  END um_iw[160]
  PIN um_iw[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 776.790 0.000 777.090 1.000 ;
    END
  END um_iw[161]
  PIN um_iw[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 839.350 53.400 839.650 54.400 ;
    END
  END um_iw[162]
  PIN um_iw[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 835.670 53.400 835.970 54.400 ;
    END
  END um_iw[163]
  PIN um_iw[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 831.990 53.400 832.290 54.400 ;
    END
  END um_iw[164]
  PIN um_iw[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 828.310 53.400 828.610 54.400 ;
    END
  END um_iw[165]
  PIN um_iw[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 824.630 53.400 824.930 54.400 ;
    END
  END um_iw[166]
  PIN um_iw[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 820.950 53.400 821.250 54.400 ;
    END
  END um_iw[167]
  PIN um_iw[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 817.270 53.400 817.570 54.400 ;
    END
  END um_iw[168]
  PIN um_iw[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 813.590 53.400 813.890 54.400 ;
    END
  END um_iw[169]
  PIN um_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 99.670 0.000 99.970 1.000 ;
    END
  END um_iw[16]
  PIN um_iw[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 809.910 53.400 810.210 54.400 ;
    END
  END um_iw[170]
  PIN um_iw[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 806.230 53.400 806.530 54.400 ;
    END
  END um_iw[171]
  PIN um_iw[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 802.550 53.400 802.850 54.400 ;
    END
  END um_iw[172]
  PIN um_iw[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 798.870 53.400 799.170 54.400 ;
    END
  END um_iw[173]
  PIN um_iw[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 795.190 53.400 795.490 54.400 ;
    END
  END um_iw[174]
  PIN um_iw[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 791.510 53.400 791.810 54.400 ;
    END
  END um_iw[175]
  PIN um_iw[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 787.830 53.400 788.130 54.400 ;
    END
  END um_iw[176]
  PIN um_iw[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 784.150 53.400 784.450 54.400 ;
    END
  END um_iw[177]
  PIN um_iw[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 780.470 53.400 780.770 54.400 ;
    END
  END um_iw[178]
  PIN um_iw[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 776.790 53.400 777.090 54.400 ;
    END
  END um_iw[179]
  PIN um_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 95.990 0.000 96.290 1.000 ;
    END
  END um_iw[17]
  PIN um_iw[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1009.550 0.000 1009.850 1.000 ;
    END
  END um_iw[180]
  PIN um_iw[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1005.870 0.000 1006.170 1.000 ;
    END
  END um_iw[181]
  PIN um_iw[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1002.190 0.000 1002.490 1.000 ;
    END
  END um_iw[182]
  PIN um_iw[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 998.510 0.000 998.810 1.000 ;
    END
  END um_iw[183]
  PIN um_iw[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 994.830 0.000 995.130 1.000 ;
    END
  END um_iw[184]
  PIN um_iw[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 991.150 0.000 991.450 1.000 ;
    END
  END um_iw[185]
  PIN um_iw[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 987.470 0.000 987.770 1.000 ;
    END
  END um_iw[186]
  PIN um_iw[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 983.790 0.000 984.090 1.000 ;
    END
  END um_iw[187]
  PIN um_iw[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 980.110 0.000 980.410 1.000 ;
    END
  END um_iw[188]
  PIN um_iw[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 976.430 0.000 976.730 1.000 ;
    END
  END um_iw[189]
  PIN um_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 158.550 53.400 158.850 54.400 ;
    END
  END um_iw[18]
  PIN um_iw[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 972.750 0.000 973.050 1.000 ;
    END
  END um_iw[190]
  PIN um_iw[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 969.070 0.000 969.370 1.000 ;
    END
  END um_iw[191]
  PIN um_iw[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 965.390 0.000 965.690 1.000 ;
    END
  END um_iw[192]
  PIN um_iw[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 961.710 0.000 962.010 1.000 ;
    END
  END um_iw[193]
  PIN um_iw[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 958.030 0.000 958.330 1.000 ;
    END
  END um_iw[194]
  PIN um_iw[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 954.350 0.000 954.650 1.000 ;
    END
  END um_iw[195]
  PIN um_iw[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 950.670 0.000 950.970 1.000 ;
    END
  END um_iw[196]
  PIN um_iw[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 946.990 0.000 947.290 1.000 ;
    END
  END um_iw[197]
  PIN um_iw[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1009.550 53.400 1009.850 54.400 ;
    END
  END um_iw[198]
  PIN um_iw[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1005.870 53.400 1006.170 54.400 ;
    END
  END um_iw[199]
  PIN um_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 154.870 53.400 155.170 54.400 ;
    END
  END um_iw[19]
  PIN um_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 154.870 0.000 155.170 1.000 ;
    END
  END um_iw[1]
  PIN um_iw[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1002.190 53.400 1002.490 54.400 ;
    END
  END um_iw[200]
  PIN um_iw[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 998.510 53.400 998.810 54.400 ;
    END
  END um_iw[201]
  PIN um_iw[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 994.830 53.400 995.130 54.400 ;
    END
  END um_iw[202]
  PIN um_iw[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 991.150 53.400 991.450 54.400 ;
    END
  END um_iw[203]
  PIN um_iw[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 987.470 53.400 987.770 54.400 ;
    END
  END um_iw[204]
  PIN um_iw[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 983.790 53.400 984.090 54.400 ;
    END
  END um_iw[205]
  PIN um_iw[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 980.110 53.400 980.410 54.400 ;
    END
  END um_iw[206]
  PIN um_iw[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 976.430 53.400 976.730 54.400 ;
    END
  END um_iw[207]
  PIN um_iw[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 972.750 53.400 973.050 54.400 ;
    END
  END um_iw[208]
  PIN um_iw[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 969.070 53.400 969.370 54.400 ;
    END
  END um_iw[209]
  PIN um_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 53.400 151.490 54.400 ;
    END
  END um_iw[20]
  PIN um_iw[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 965.390 53.400 965.690 54.400 ;
    END
  END um_iw[210]
  PIN um_iw[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 961.710 53.400 962.010 54.400 ;
    END
  END um_iw[211]
  PIN um_iw[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 958.030 53.400 958.330 54.400 ;
    END
  END um_iw[212]
  PIN um_iw[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 954.350 53.400 954.650 54.400 ;
    END
  END um_iw[213]
  PIN um_iw[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 950.670 53.400 950.970 54.400 ;
    END
  END um_iw[214]
  PIN um_iw[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 946.990 53.400 947.290 54.400 ;
    END
  END um_iw[215]
  PIN um_iw[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1179.750 0.000 1180.050 1.000 ;
    END
  END um_iw[216]
  PIN um_iw[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1176.070 0.000 1176.370 1.000 ;
    END
  END um_iw[217]
  PIN um_iw[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1172.390 0.000 1172.690 1.000 ;
    END
  END um_iw[218]
  PIN um_iw[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1168.710 0.000 1169.010 1.000 ;
    END
  END um_iw[219]
  PIN um_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 53.400 147.810 54.400 ;
    END
  END um_iw[21]
  PIN um_iw[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1165.030 0.000 1165.330 1.000 ;
    END
  END um_iw[220]
  PIN um_iw[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1161.350 0.000 1161.650 1.000 ;
    END
  END um_iw[221]
  PIN um_iw[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1157.670 0.000 1157.970 1.000 ;
    END
  END um_iw[222]
  PIN um_iw[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1153.990 0.000 1154.290 1.000 ;
    END
  END um_iw[223]
  PIN um_iw[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1150.310 0.000 1150.610 1.000 ;
    END
  END um_iw[224]
  PIN um_iw[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1146.630 0.000 1146.930 1.000 ;
    END
  END um_iw[225]
  PIN um_iw[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1142.950 0.000 1143.250 1.000 ;
    END
  END um_iw[226]
  PIN um_iw[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1139.270 0.000 1139.570 1.000 ;
    END
  END um_iw[227]
  PIN um_iw[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1135.590 0.000 1135.890 1.000 ;
    END
  END um_iw[228]
  PIN um_iw[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1131.910 0.000 1132.210 1.000 ;
    END
  END um_iw[229]
  PIN um_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 53.400 144.130 54.400 ;
    END
  END um_iw[22]
  PIN um_iw[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1128.230 0.000 1128.530 1.000 ;
    END
  END um_iw[230]
  PIN um_iw[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1124.550 0.000 1124.850 1.000 ;
    END
  END um_iw[231]
  PIN um_iw[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1120.870 0.000 1121.170 1.000 ;
    END
  END um_iw[232]
  PIN um_iw[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1117.190 0.000 1117.490 1.000 ;
    END
  END um_iw[233]
  PIN um_iw[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1179.750 53.400 1180.050 54.400 ;
    END
  END um_iw[234]
  PIN um_iw[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1176.070 53.400 1176.370 54.400 ;
    END
  END um_iw[235]
  PIN um_iw[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1172.390 53.400 1172.690 54.400 ;
    END
  END um_iw[236]
  PIN um_iw[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1168.710 53.400 1169.010 54.400 ;
    END
  END um_iw[237]
  PIN um_iw[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1165.030 53.400 1165.330 54.400 ;
    END
  END um_iw[238]
  PIN um_iw[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1161.350 53.400 1161.650 54.400 ;
    END
  END um_iw[239]
  PIN um_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 53.400 140.450 54.400 ;
    END
  END um_iw[23]
  PIN um_iw[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1157.670 53.400 1157.970 54.400 ;
    END
  END um_iw[240]
  PIN um_iw[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1153.990 53.400 1154.290 54.400 ;
    END
  END um_iw[241]
  PIN um_iw[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1150.310 53.400 1150.610 54.400 ;
    END
  END um_iw[242]
  PIN um_iw[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1146.630 53.400 1146.930 54.400 ;
    END
  END um_iw[243]
  PIN um_iw[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1142.950 53.400 1143.250 54.400 ;
    END
  END um_iw[244]
  PIN um_iw[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1139.270 53.400 1139.570 54.400 ;
    END
  END um_iw[245]
  PIN um_iw[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1135.590 53.400 1135.890 54.400 ;
    END
  END um_iw[246]
  PIN um_iw[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1131.910 53.400 1132.210 54.400 ;
    END
  END um_iw[247]
  PIN um_iw[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1128.230 53.400 1128.530 54.400 ;
    END
  END um_iw[248]
  PIN um_iw[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1124.550 53.400 1124.850 54.400 ;
    END
  END um_iw[249]
  PIN um_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 53.400 136.770 54.400 ;
    END
  END um_iw[24]
  PIN um_iw[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1120.870 53.400 1121.170 54.400 ;
    END
  END um_iw[250]
  PIN um_iw[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1117.190 53.400 1117.490 54.400 ;
    END
  END um_iw[251]
  PIN um_iw[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1349.950 0.000 1350.250 1.000 ;
    END
  END um_iw[252]
  PIN um_iw[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1346.270 0.000 1346.570 1.000 ;
    END
  END um_iw[253]
  PIN um_iw[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1342.590 0.000 1342.890 1.000 ;
    END
  END um_iw[254]
  PIN um_iw[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1338.910 0.000 1339.210 1.000 ;
    END
  END um_iw[255]
  PIN um_iw[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1335.230 0.000 1335.530 1.000 ;
    END
  END um_iw[256]
  PIN um_iw[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1331.550 0.000 1331.850 1.000 ;
    END
  END um_iw[257]
  PIN um_iw[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1327.870 0.000 1328.170 1.000 ;
    END
  END um_iw[258]
  PIN um_iw[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1324.190 0.000 1324.490 1.000 ;
    END
  END um_iw[259]
  PIN um_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 53.400 133.090 54.400 ;
    END
  END um_iw[25]
  PIN um_iw[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1320.510 0.000 1320.810 1.000 ;
    END
  END um_iw[260]
  PIN um_iw[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1316.830 0.000 1317.130 1.000 ;
    END
  END um_iw[261]
  PIN um_iw[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1313.150 0.000 1313.450 1.000 ;
    END
  END um_iw[262]
  PIN um_iw[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1309.470 0.000 1309.770 1.000 ;
    END
  END um_iw[263]
  PIN um_iw[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1305.790 0.000 1306.090 1.000 ;
    END
  END um_iw[264]
  PIN um_iw[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1302.110 0.000 1302.410 1.000 ;
    END
  END um_iw[265]
  PIN um_iw[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1298.430 0.000 1298.730 1.000 ;
    END
  END um_iw[266]
  PIN um_iw[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1294.750 0.000 1295.050 1.000 ;
    END
  END um_iw[267]
  PIN um_iw[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1291.070 0.000 1291.370 1.000 ;
    END
  END um_iw[268]
  PIN um_iw[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1287.390 0.000 1287.690 1.000 ;
    END
  END um_iw[269]
  PIN um_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 53.400 129.410 54.400 ;
    END
  END um_iw[26]
  PIN um_iw[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1349.950 53.400 1350.250 54.400 ;
    END
  END um_iw[270]
  PIN um_iw[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1346.270 53.400 1346.570 54.400 ;
    END
  END um_iw[271]
  PIN um_iw[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1342.590 53.400 1342.890 54.400 ;
    END
  END um_iw[272]
  PIN um_iw[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1338.910 53.400 1339.210 54.400 ;
    END
  END um_iw[273]
  PIN um_iw[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1335.230 53.400 1335.530 54.400 ;
    END
  END um_iw[274]
  PIN um_iw[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1331.550 53.400 1331.850 54.400 ;
    END
  END um_iw[275]
  PIN um_iw[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1327.870 53.400 1328.170 54.400 ;
    END
  END um_iw[276]
  PIN um_iw[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1324.190 53.400 1324.490 54.400 ;
    END
  END um_iw[277]
  PIN um_iw[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1320.510 53.400 1320.810 54.400 ;
    END
  END um_iw[278]
  PIN um_iw[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1316.830 53.400 1317.130 54.400 ;
    END
  END um_iw[279]
  PIN um_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 53.400 125.730 54.400 ;
    END
  END um_iw[27]
  PIN um_iw[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1313.150 53.400 1313.450 54.400 ;
    END
  END um_iw[280]
  PIN um_iw[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1309.470 53.400 1309.770 54.400 ;
    END
  END um_iw[281]
  PIN um_iw[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1305.790 53.400 1306.090 54.400 ;
    END
  END um_iw[282]
  PIN um_iw[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1302.110 53.400 1302.410 54.400 ;
    END
  END um_iw[283]
  PIN um_iw[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1298.430 53.400 1298.730 54.400 ;
    END
  END um_iw[284]
  PIN um_iw[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1294.750 53.400 1295.050 54.400 ;
    END
  END um_iw[285]
  PIN um_iw[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1291.070 53.400 1291.370 54.400 ;
    END
  END um_iw[286]
  PIN um_iw[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1287.390 53.400 1287.690 54.400 ;
    END
  END um_iw[287]
  PIN um_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 53.400 122.050 54.400 ;
    END
  END um_iw[28]
  PIN um_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 53.400 118.370 54.400 ;
    END
  END um_iw[29]
  PIN um_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 0.000 151.490 1.000 ;
    END
  END um_iw[2]
  PIN um_iw[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 53.400 114.690 54.400 ;
    END
  END um_iw[30]
  PIN um_iw[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 53.400 111.010 54.400 ;
    END
  END um_iw[31]
  PIN um_iw[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 53.400 107.330 54.400 ;
    END
  END um_iw[32]
  PIN um_iw[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 103.350 53.400 103.650 54.400 ;
    END
  END um_iw[33]
  PIN um_iw[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 99.670 53.400 99.970 54.400 ;
    END
  END um_iw[34]
  PIN um_iw[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 95.990 53.400 96.290 54.400 ;
    END
  END um_iw[35]
  PIN um_iw[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 328.750 0.000 329.050 1.000 ;
    END
  END um_iw[36]
  PIN um_iw[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 325.070 0.000 325.370 1.000 ;
    END
  END um_iw[37]
  PIN um_iw[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 321.390 0.000 321.690 1.000 ;
    END
  END um_iw[38]
  PIN um_iw[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 317.710 0.000 318.010 1.000 ;
    END
  END um_iw[39]
  PIN um_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 0.000 147.810 1.000 ;
    END
  END um_iw[3]
  PIN um_iw[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 314.030 0.000 314.330 1.000 ;
    END
  END um_iw[40]
  PIN um_iw[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 310.350 0.000 310.650 1.000 ;
    END
  END um_iw[41]
  PIN um_iw[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 306.670 0.000 306.970 1.000 ;
    END
  END um_iw[42]
  PIN um_iw[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 302.990 0.000 303.290 1.000 ;
    END
  END um_iw[43]
  PIN um_iw[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 299.310 0.000 299.610 1.000 ;
    END
  END um_iw[44]
  PIN um_iw[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 295.630 0.000 295.930 1.000 ;
    END
  END um_iw[45]
  PIN um_iw[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 291.950 0.000 292.250 1.000 ;
    END
  END um_iw[46]
  PIN um_iw[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 288.270 0.000 288.570 1.000 ;
    END
  END um_iw[47]
  PIN um_iw[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 284.590 0.000 284.890 1.000 ;
    END
  END um_iw[48]
  PIN um_iw[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 280.910 0.000 281.210 1.000 ;
    END
  END um_iw[49]
  PIN um_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 0.000 144.130 1.000 ;
    END
  END um_iw[4]
  PIN um_iw[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 277.230 0.000 277.530 1.000 ;
    END
  END um_iw[50]
  PIN um_iw[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 273.550 0.000 273.850 1.000 ;
    END
  END um_iw[51]
  PIN um_iw[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 269.870 0.000 270.170 1.000 ;
    END
  END um_iw[52]
  PIN um_iw[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 266.190 0.000 266.490 1.000 ;
    END
  END um_iw[53]
  PIN um_iw[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 328.750 53.400 329.050 54.400 ;
    END
  END um_iw[54]
  PIN um_iw[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 325.070 53.400 325.370 54.400 ;
    END
  END um_iw[55]
  PIN um_iw[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 321.390 53.400 321.690 54.400 ;
    END
  END um_iw[56]
  PIN um_iw[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 317.710 53.400 318.010 54.400 ;
    END
  END um_iw[57]
  PIN um_iw[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 314.030 53.400 314.330 54.400 ;
    END
  END um_iw[58]
  PIN um_iw[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 310.350 53.400 310.650 54.400 ;
    END
  END um_iw[59]
  PIN um_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 0.000 140.450 1.000 ;
    END
  END um_iw[5]
  PIN um_iw[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 306.670 53.400 306.970 54.400 ;
    END
  END um_iw[60]
  PIN um_iw[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 302.990 53.400 303.290 54.400 ;
    END
  END um_iw[61]
  PIN um_iw[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 299.310 53.400 299.610 54.400 ;
    END
  END um_iw[62]
  PIN um_iw[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 295.630 53.400 295.930 54.400 ;
    END
  END um_iw[63]
  PIN um_iw[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 291.950 53.400 292.250 54.400 ;
    END
  END um_iw[64]
  PIN um_iw[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 288.270 53.400 288.570 54.400 ;
    END
  END um_iw[65]
  PIN um_iw[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 284.590 53.400 284.890 54.400 ;
    END
  END um_iw[66]
  PIN um_iw[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 280.910 53.400 281.210 54.400 ;
    END
  END um_iw[67]
  PIN um_iw[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 277.230 53.400 277.530 54.400 ;
    END
  END um_iw[68]
  PIN um_iw[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 273.550 53.400 273.850 54.400 ;
    END
  END um_iw[69]
  PIN um_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 0.000 136.770 1.000 ;
    END
  END um_iw[6]
  PIN um_iw[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 269.870 53.400 270.170 54.400 ;
    END
  END um_iw[70]
  PIN um_iw[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 266.190 53.400 266.490 54.400 ;
    END
  END um_iw[71]
  PIN um_iw[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 498.950 0.000 499.250 1.000 ;
    END
  END um_iw[72]
  PIN um_iw[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 495.270 0.000 495.570 1.000 ;
    END
  END um_iw[73]
  PIN um_iw[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 491.590 0.000 491.890 1.000 ;
    END
  END um_iw[74]
  PIN um_iw[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 487.910 0.000 488.210 1.000 ;
    END
  END um_iw[75]
  PIN um_iw[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 484.230 0.000 484.530 1.000 ;
    END
  END um_iw[76]
  PIN um_iw[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 480.550 0.000 480.850 1.000 ;
    END
  END um_iw[77]
  PIN um_iw[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 476.870 0.000 477.170 1.000 ;
    END
  END um_iw[78]
  PIN um_iw[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 473.190 0.000 473.490 1.000 ;
    END
  END um_iw[79]
  PIN um_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 0.000 133.090 1.000 ;
    END
  END um_iw[7]
  PIN um_iw[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 469.510 0.000 469.810 1.000 ;
    END
  END um_iw[80]
  PIN um_iw[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 465.830 0.000 466.130 1.000 ;
    END
  END um_iw[81]
  PIN um_iw[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 462.150 0.000 462.450 1.000 ;
    END
  END um_iw[82]
  PIN um_iw[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 458.470 0.000 458.770 1.000 ;
    END
  END um_iw[83]
  PIN um_iw[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 454.790 0.000 455.090 1.000 ;
    END
  END um_iw[84]
  PIN um_iw[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 451.110 0.000 451.410 1.000 ;
    END
  END um_iw[85]
  PIN um_iw[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 447.430 0.000 447.730 1.000 ;
    END
  END um_iw[86]
  PIN um_iw[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 443.750 0.000 444.050 1.000 ;
    END
  END um_iw[87]
  PIN um_iw[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 440.070 0.000 440.370 1.000 ;
    END
  END um_iw[88]
  PIN um_iw[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 436.390 0.000 436.690 1.000 ;
    END
  END um_iw[89]
  PIN um_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 0.000 129.410 1.000 ;
    END
  END um_iw[8]
  PIN um_iw[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 498.950 53.400 499.250 54.400 ;
    END
  END um_iw[90]
  PIN um_iw[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 495.270 53.400 495.570 54.400 ;
    END
  END um_iw[91]
  PIN um_iw[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 491.590 53.400 491.890 54.400 ;
    END
  END um_iw[92]
  PIN um_iw[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 487.910 53.400 488.210 54.400 ;
    END
  END um_iw[93]
  PIN um_iw[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 484.230 53.400 484.530 54.400 ;
    END
  END um_iw[94]
  PIN um_iw[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 480.550 53.400 480.850 54.400 ;
    END
  END um_iw[95]
  PIN um_iw[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 476.870 53.400 477.170 54.400 ;
    END
  END um_iw[96]
  PIN um_iw[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 473.190 53.400 473.490 54.400 ;
    END
  END um_iw[97]
  PIN um_iw[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 469.510 53.400 469.810 54.400 ;
    END
  END um_iw[98]
  PIN um_iw[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 465.830 53.400 466.130 54.400 ;
    END
  END um_iw[99]
  PIN um_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 0.000 125.730 1.000 ;
    END
  END um_iw[9]
  PIN um_k_zero[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 0.000 4.290 1.000 ;
    END
  END um_k_zero[0]
  PIN um_k_zero[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 854.990 0.000 855.290 1.000 ;
    END
  END um_k_zero[10]
  PIN um_k_zero[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 854.990 53.400 855.290 54.400 ;
    END
  END um_k_zero[11]
  PIN um_k_zero[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1025.190 0.000 1025.490 1.000 ;
    END
  END um_k_zero[12]
  PIN um_k_zero[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1025.190 53.400 1025.490 54.400 ;
    END
  END um_k_zero[13]
  PIN um_k_zero[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1195.390 0.000 1195.690 1.000 ;
    END
  END um_k_zero[14]
  PIN um_k_zero[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1195.390 53.400 1195.690 54.400 ;
    END
  END um_k_zero[15]
  PIN um_k_zero[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 53.400 4.290 54.400 ;
    END
  END um_k_zero[1]
  PIN um_k_zero[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 174.190 0.000 174.490 1.000 ;
    END
  END um_k_zero[2]
  PIN um_k_zero[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 174.190 53.400 174.490 54.400 ;
    END
  END um_k_zero[3]
  PIN um_k_zero[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 344.390 0.000 344.690 1.000 ;
    END
  END um_k_zero[4]
  PIN um_k_zero[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 344.390 53.400 344.690 54.400 ;
    END
  END um_k_zero[5]
  PIN um_k_zero[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 514.590 0.000 514.890 1.000 ;
    END
  END um_k_zero[6]
  PIN um_k_zero[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 514.590 53.400 514.890 54.400 ;
    END
  END um_k_zero[7]
  PIN um_k_zero[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 684.790 0.000 685.090 1.000 ;
    END
  END um_k_zero[8]
  PIN um_k_zero[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 684.790 53.400 685.090 54.400 ;
    END
  END um_k_zero[9]
  PIN um_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 0.000 92.610 1.000 ;
    END
  END um_ow[0]
  PIN um_ow[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 417.990 0.000 418.290 1.000 ;
    END
  END um_ow[100]
  PIN um_ow[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 414.310 0.000 414.610 1.000 ;
    END
  END um_ow[101]
  PIN um_ow[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 410.630 0.000 410.930 1.000 ;
    END
  END um_ow[102]
  PIN um_ow[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 406.950 0.000 407.250 1.000 ;
    END
  END um_ow[103]
  PIN um_ow[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 403.270 0.000 403.570 1.000 ;
    END
  END um_ow[104]
  PIN um_ow[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 399.590 0.000 399.890 1.000 ;
    END
  END um_ow[105]
  PIN um_ow[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 395.910 0.000 396.210 1.000 ;
    END
  END um_ow[106]
  PIN um_ow[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 392.230 0.000 392.530 1.000 ;
    END
  END um_ow[107]
  PIN um_ow[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 388.550 0.000 388.850 1.000 ;
    END
  END um_ow[108]
  PIN um_ow[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 384.870 0.000 385.170 1.000 ;
    END
  END um_ow[109]
  PIN um_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 55.510 0.000 55.810 1.000 ;
    END
  END um_ow[10]
  PIN um_ow[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 381.190 0.000 381.490 1.000 ;
    END
  END um_ow[110]
  PIN um_ow[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 377.510 0.000 377.810 1.000 ;
    END
  END um_ow[111]
  PIN um_ow[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 373.830 0.000 374.130 1.000 ;
    END
  END um_ow[112]
  PIN um_ow[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 370.150 0.000 370.450 1.000 ;
    END
  END um_ow[113]
  PIN um_ow[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 366.470 0.000 366.770 1.000 ;
    END
  END um_ow[114]
  PIN um_ow[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 362.790 0.000 363.090 1.000 ;
    END
  END um_ow[115]
  PIN um_ow[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 359.110 0.000 359.410 1.000 ;
    END
  END um_ow[116]
  PIN um_ow[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 355.430 0.000 355.730 1.000 ;
    END
  END um_ow[117]
  PIN um_ow[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 351.750 0.000 352.050 1.000 ;
    END
  END um_ow[118]
  PIN um_ow[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 348.070 0.000 348.370 1.000 ;
    END
  END um_ow[119]
  PIN um_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 51.830 0.000 52.130 1.000 ;
    END
  END um_ow[11]
  PIN um_ow[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 432.710 53.400 433.010 54.400 ;
    END
  END um_ow[120]
  PIN um_ow[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 429.030 53.400 429.330 54.400 ;
    END
  END um_ow[121]
  PIN um_ow[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 425.350 53.400 425.650 54.400 ;
    END
  END um_ow[122]
  PIN um_ow[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 421.670 53.400 421.970 54.400 ;
    END
  END um_ow[123]
  PIN um_ow[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 417.990 53.400 418.290 54.400 ;
    END
  END um_ow[124]
  PIN um_ow[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 414.310 53.400 414.610 54.400 ;
    END
  END um_ow[125]
  PIN um_ow[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 410.630 53.400 410.930 54.400 ;
    END
  END um_ow[126]
  PIN um_ow[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 406.950 53.400 407.250 54.400 ;
    END
  END um_ow[127]
  PIN um_ow[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 403.270 53.400 403.570 54.400 ;
    END
  END um_ow[128]
  PIN um_ow[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 399.590 53.400 399.890 54.400 ;
    END
  END um_ow[129]
  PIN um_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 48.150 0.000 48.450 1.000 ;
    END
  END um_ow[12]
  PIN um_ow[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 395.910 53.400 396.210 54.400 ;
    END
  END um_ow[130]
  PIN um_ow[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 392.230 53.400 392.530 54.400 ;
    END
  END um_ow[131]
  PIN um_ow[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 388.550 53.400 388.850 54.400 ;
    END
  END um_ow[132]
  PIN um_ow[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 384.870 53.400 385.170 54.400 ;
    END
  END um_ow[133]
  PIN um_ow[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 381.190 53.400 381.490 54.400 ;
    END
  END um_ow[134]
  PIN um_ow[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 377.510 53.400 377.810 54.400 ;
    END
  END um_ow[135]
  PIN um_ow[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 373.830 53.400 374.130 54.400 ;
    END
  END um_ow[136]
  PIN um_ow[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 370.150 53.400 370.450 54.400 ;
    END
  END um_ow[137]
  PIN um_ow[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 366.470 53.400 366.770 54.400 ;
    END
  END um_ow[138]
  PIN um_ow[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 362.790 53.400 363.090 54.400 ;
    END
  END um_ow[139]
  PIN um_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 0.000 44.770 1.000 ;
    END
  END um_ow[13]
  PIN um_ow[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 359.110 53.400 359.410 54.400 ;
    END
  END um_ow[140]
  PIN um_ow[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 355.430 53.400 355.730 54.400 ;
    END
  END um_ow[141]
  PIN um_ow[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 351.750 53.400 352.050 54.400 ;
    END
  END um_ow[142]
  PIN um_ow[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 348.070 53.400 348.370 54.400 ;
    END
  END um_ow[143]
  PIN um_ow[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 602.910 0.000 603.210 1.000 ;
    END
  END um_ow[144]
  PIN um_ow[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 599.230 0.000 599.530 1.000 ;
    END
  END um_ow[145]
  PIN um_ow[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 595.550 0.000 595.850 1.000 ;
    END
  END um_ow[146]
  PIN um_ow[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 591.870 0.000 592.170 1.000 ;
    END
  END um_ow[147]
  PIN um_ow[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 588.190 0.000 588.490 1.000 ;
    END
  END um_ow[148]
  PIN um_ow[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 584.510 0.000 584.810 1.000 ;
    END
  END um_ow[149]
  PIN um_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 0.000 41.090 1.000 ;
    END
  END um_ow[14]
  PIN um_ow[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 580.830 0.000 581.130 1.000 ;
    END
  END um_ow[150]
  PIN um_ow[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 577.150 0.000 577.450 1.000 ;
    END
  END um_ow[151]
  PIN um_ow[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 573.470 0.000 573.770 1.000 ;
    END
  END um_ow[152]
  PIN um_ow[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 569.790 0.000 570.090 1.000 ;
    END
  END um_ow[153]
  PIN um_ow[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 566.110 0.000 566.410 1.000 ;
    END
  END um_ow[154]
  PIN um_ow[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 562.430 0.000 562.730 1.000 ;
    END
  END um_ow[155]
  PIN um_ow[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 558.750 0.000 559.050 1.000 ;
    END
  END um_ow[156]
  PIN um_ow[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 555.070 0.000 555.370 1.000 ;
    END
  END um_ow[157]
  PIN um_ow[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 551.390 0.000 551.690 1.000 ;
    END
  END um_ow[158]
  PIN um_ow[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 547.710 0.000 548.010 1.000 ;
    END
  END um_ow[159]
  PIN um_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 37.110 0.000 37.410 1.000 ;
    END
  END um_ow[15]
  PIN um_ow[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 544.030 0.000 544.330 1.000 ;
    END
  END um_ow[160]
  PIN um_ow[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 540.350 0.000 540.650 1.000 ;
    END
  END um_ow[161]
  PIN um_ow[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 536.670 0.000 536.970 1.000 ;
    END
  END um_ow[162]
  PIN um_ow[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 532.990 0.000 533.290 1.000 ;
    END
  END um_ow[163]
  PIN um_ow[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 529.310 0.000 529.610 1.000 ;
    END
  END um_ow[164]
  PIN um_ow[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 525.630 0.000 525.930 1.000 ;
    END
  END um_ow[165]
  PIN um_ow[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 521.950 0.000 522.250 1.000 ;
    END
  END um_ow[166]
  PIN um_ow[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 518.270 0.000 518.570 1.000 ;
    END
  END um_ow[167]
  PIN um_ow[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 602.910 53.400 603.210 54.400 ;
    END
  END um_ow[168]
  PIN um_ow[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 599.230 53.400 599.530 54.400 ;
    END
  END um_ow[169]
  PIN um_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 33.430 0.000 33.730 1.000 ;
    END
  END um_ow[16]
  PIN um_ow[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 595.550 53.400 595.850 54.400 ;
    END
  END um_ow[170]
  PIN um_ow[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 591.870 53.400 592.170 54.400 ;
    END
  END um_ow[171]
  PIN um_ow[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 588.190 53.400 588.490 54.400 ;
    END
  END um_ow[172]
  PIN um_ow[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 584.510 53.400 584.810 54.400 ;
    END
  END um_ow[173]
  PIN um_ow[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 580.830 53.400 581.130 54.400 ;
    END
  END um_ow[174]
  PIN um_ow[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 577.150 53.400 577.450 54.400 ;
    END
  END um_ow[175]
  PIN um_ow[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 573.470 53.400 573.770 54.400 ;
    END
  END um_ow[176]
  PIN um_ow[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 569.790 53.400 570.090 54.400 ;
    END
  END um_ow[177]
  PIN um_ow[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 566.110 53.400 566.410 54.400 ;
    END
  END um_ow[178]
  PIN um_ow[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 562.430 53.400 562.730 54.400 ;
    END
  END um_ow[179]
  PIN um_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 29.750 0.000 30.050 1.000 ;
    END
  END um_ow[17]
  PIN um_ow[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 558.750 53.400 559.050 54.400 ;
    END
  END um_ow[180]
  PIN um_ow[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 555.070 53.400 555.370 54.400 ;
    END
  END um_ow[181]
  PIN um_ow[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 551.390 53.400 551.690 54.400 ;
    END
  END um_ow[182]
  PIN um_ow[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 547.710 53.400 548.010 54.400 ;
    END
  END um_ow[183]
  PIN um_ow[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 544.030 53.400 544.330 54.400 ;
    END
  END um_ow[184]
  PIN um_ow[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 540.350 53.400 540.650 54.400 ;
    END
  END um_ow[185]
  PIN um_ow[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 536.670 53.400 536.970 54.400 ;
    END
  END um_ow[186]
  PIN um_ow[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 532.990 53.400 533.290 54.400 ;
    END
  END um_ow[187]
  PIN um_ow[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 529.310 53.400 529.610 54.400 ;
    END
  END um_ow[188]
  PIN um_ow[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 525.630 53.400 525.930 54.400 ;
    END
  END um_ow[189]
  PIN um_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 26.070 0.000 26.370 1.000 ;
    END
  END um_ow[18]
  PIN um_ow[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 521.950 53.400 522.250 54.400 ;
    END
  END um_ow[190]
  PIN um_ow[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 518.270 53.400 518.570 54.400 ;
    END
  END um_ow[191]
  PIN um_ow[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 773.110 0.000 773.410 1.000 ;
    END
  END um_ow[192]
  PIN um_ow[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 769.430 0.000 769.730 1.000 ;
    END
  END um_ow[193]
  PIN um_ow[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 765.750 0.000 766.050 1.000 ;
    END
  END um_ow[194]
  PIN um_ow[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 762.070 0.000 762.370 1.000 ;
    END
  END um_ow[195]
  PIN um_ow[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 758.390 0.000 758.690 1.000 ;
    END
  END um_ow[196]
  PIN um_ow[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 754.710 0.000 755.010 1.000 ;
    END
  END um_ow[197]
  PIN um_ow[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 751.030 0.000 751.330 1.000 ;
    END
  END um_ow[198]
  PIN um_ow[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 747.350 0.000 747.650 1.000 ;
    END
  END um_ow[199]
  PIN um_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 22.390 0.000 22.690 1.000 ;
    END
  END um_ow[19]
  PIN um_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 88.630 0.000 88.930 1.000 ;
    END
  END um_ow[1]
  PIN um_ow[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 743.670 0.000 743.970 1.000 ;
    END
  END um_ow[200]
  PIN um_ow[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 739.990 0.000 740.290 1.000 ;
    END
  END um_ow[201]
  PIN um_ow[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 736.310 0.000 736.610 1.000 ;
    END
  END um_ow[202]
  PIN um_ow[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 732.630 0.000 732.930 1.000 ;
    END
  END um_ow[203]
  PIN um_ow[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 728.950 0.000 729.250 1.000 ;
    END
  END um_ow[204]
  PIN um_ow[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 725.270 0.000 725.570 1.000 ;
    END
  END um_ow[205]
  PIN um_ow[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 721.590 0.000 721.890 1.000 ;
    END
  END um_ow[206]
  PIN um_ow[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 717.910 0.000 718.210 1.000 ;
    END
  END um_ow[207]
  PIN um_ow[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 714.230 0.000 714.530 1.000 ;
    END
  END um_ow[208]
  PIN um_ow[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 710.550 0.000 710.850 1.000 ;
    END
  END um_ow[209]
  PIN um_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 18.710 0.000 19.010 1.000 ;
    END
  END um_ow[20]
  PIN um_ow[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 706.870 0.000 707.170 1.000 ;
    END
  END um_ow[210]
  PIN um_ow[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 703.190 0.000 703.490 1.000 ;
    END
  END um_ow[211]
  PIN um_ow[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 699.510 0.000 699.810 1.000 ;
    END
  END um_ow[212]
  PIN um_ow[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 695.830 0.000 696.130 1.000 ;
    END
  END um_ow[213]
  PIN um_ow[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 692.150 0.000 692.450 1.000 ;
    END
  END um_ow[214]
  PIN um_ow[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 688.470 0.000 688.770 1.000 ;
    END
  END um_ow[215]
  PIN um_ow[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 773.110 53.400 773.410 54.400 ;
    END
  END um_ow[216]
  PIN um_ow[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 769.430 53.400 769.730 54.400 ;
    END
  END um_ow[217]
  PIN um_ow[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 765.750 53.400 766.050 54.400 ;
    END
  END um_ow[218]
  PIN um_ow[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 762.070 53.400 762.370 54.400 ;
    END
  END um_ow[219]
  PIN um_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 15.030 0.000 15.330 1.000 ;
    END
  END um_ow[21]
  PIN um_ow[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 758.390 53.400 758.690 54.400 ;
    END
  END um_ow[220]
  PIN um_ow[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 754.710 53.400 755.010 54.400 ;
    END
  END um_ow[221]
  PIN um_ow[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 751.030 53.400 751.330 54.400 ;
    END
  END um_ow[222]
  PIN um_ow[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 747.350 53.400 747.650 54.400 ;
    END
  END um_ow[223]
  PIN um_ow[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 743.670 53.400 743.970 54.400 ;
    END
  END um_ow[224]
  PIN um_ow[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 739.990 53.400 740.290 54.400 ;
    END
  END um_ow[225]
  PIN um_ow[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 736.310 53.400 736.610 54.400 ;
    END
  END um_ow[226]
  PIN um_ow[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 732.630 53.400 732.930 54.400 ;
    END
  END um_ow[227]
  PIN um_ow[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 728.950 53.400 729.250 54.400 ;
    END
  END um_ow[228]
  PIN um_ow[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 725.270 53.400 725.570 54.400 ;
    END
  END um_ow[229]
  PIN um_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 11.350 0.000 11.650 1.000 ;
    END
  END um_ow[22]
  PIN um_ow[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 721.590 53.400 721.890 54.400 ;
    END
  END um_ow[230]
  PIN um_ow[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 717.910 53.400 718.210 54.400 ;
    END
  END um_ow[231]
  PIN um_ow[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 714.230 53.400 714.530 54.400 ;
    END
  END um_ow[232]
  PIN um_ow[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 710.550 53.400 710.850 54.400 ;
    END
  END um_ow[233]
  PIN um_ow[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 706.870 53.400 707.170 54.400 ;
    END
  END um_ow[234]
  PIN um_ow[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 703.190 53.400 703.490 54.400 ;
    END
  END um_ow[235]
  PIN um_ow[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 699.510 53.400 699.810 54.400 ;
    END
  END um_ow[236]
  PIN um_ow[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 695.830 53.400 696.130 54.400 ;
    END
  END um_ow[237]
  PIN um_ow[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 692.150 53.400 692.450 54.400 ;
    END
  END um_ow[238]
  PIN um_ow[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 688.470 53.400 688.770 54.400 ;
    END
  END um_ow[239]
  PIN um_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 7.670 0.000 7.970 1.000 ;
    END
  END um_ow[23]
  PIN um_ow[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 943.310 0.000 943.610 1.000 ;
    END
  END um_ow[240]
  PIN um_ow[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 939.630 0.000 939.930 1.000 ;
    END
  END um_ow[241]
  PIN um_ow[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 935.950 0.000 936.250 1.000 ;
    END
  END um_ow[242]
  PIN um_ow[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 932.270 0.000 932.570 1.000 ;
    END
  END um_ow[243]
  PIN um_ow[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 928.590 0.000 928.890 1.000 ;
    END
  END um_ow[244]
  PIN um_ow[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 924.910 0.000 925.210 1.000 ;
    END
  END um_ow[245]
  PIN um_ow[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 921.230 0.000 921.530 1.000 ;
    END
  END um_ow[246]
  PIN um_ow[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 917.550 0.000 917.850 1.000 ;
    END
  END um_ow[247]
  PIN um_ow[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 913.870 0.000 914.170 1.000 ;
    END
  END um_ow[248]
  PIN um_ow[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 910.190 0.000 910.490 1.000 ;
    END
  END um_ow[249]
  PIN um_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 53.400 92.610 54.400 ;
    END
  END um_ow[24]
  PIN um_ow[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 906.510 0.000 906.810 1.000 ;
    END
  END um_ow[250]
  PIN um_ow[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 902.830 0.000 903.130 1.000 ;
    END
  END um_ow[251]
  PIN um_ow[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 899.150 0.000 899.450 1.000 ;
    END
  END um_ow[252]
  PIN um_ow[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 895.470 0.000 895.770 1.000 ;
    END
  END um_ow[253]
  PIN um_ow[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 891.790 0.000 892.090 1.000 ;
    END
  END um_ow[254]
  PIN um_ow[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 888.110 0.000 888.410 1.000 ;
    END
  END um_ow[255]
  PIN um_ow[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 884.430 0.000 884.730 1.000 ;
    END
  END um_ow[256]
  PIN um_ow[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 880.750 0.000 881.050 1.000 ;
    END
  END um_ow[257]
  PIN um_ow[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 877.070 0.000 877.370 1.000 ;
    END
  END um_ow[258]
  PIN um_ow[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 873.390 0.000 873.690 1.000 ;
    END
  END um_ow[259]
  PIN um_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 53.400 88.930 54.400 ;
    END
  END um_ow[25]
  PIN um_ow[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 869.710 0.000 870.010 1.000 ;
    END
  END um_ow[260]
  PIN um_ow[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 866.030 0.000 866.330 1.000 ;
    END
  END um_ow[261]
  PIN um_ow[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 862.350 0.000 862.650 1.000 ;
    END
  END um_ow[262]
  PIN um_ow[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 858.670 0.000 858.970 1.000 ;
    END
  END um_ow[263]
  PIN um_ow[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 943.310 53.400 943.610 54.400 ;
    END
  END um_ow[264]
  PIN um_ow[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 939.630 53.400 939.930 54.400 ;
    END
  END um_ow[265]
  PIN um_ow[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 935.950 53.400 936.250 54.400 ;
    END
  END um_ow[266]
  PIN um_ow[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 932.270 53.400 932.570 54.400 ;
    END
  END um_ow[267]
  PIN um_ow[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 928.590 53.400 928.890 54.400 ;
    END
  END um_ow[268]
  PIN um_ow[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 924.910 53.400 925.210 54.400 ;
    END
  END um_ow[269]
  PIN um_ow[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.950 53.400 85.250 54.400 ;
    END
  END um_ow[26]
  PIN um_ow[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 921.230 53.400 921.530 54.400 ;
    END
  END um_ow[270]
  PIN um_ow[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 917.550 53.400 917.850 54.400 ;
    END
  END um_ow[271]
  PIN um_ow[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 913.870 53.400 914.170 54.400 ;
    END
  END um_ow[272]
  PIN um_ow[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 910.190 53.400 910.490 54.400 ;
    END
  END um_ow[273]
  PIN um_ow[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 906.510 53.400 906.810 54.400 ;
    END
  END um_ow[274]
  PIN um_ow[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 902.830 53.400 903.130 54.400 ;
    END
  END um_ow[275]
  PIN um_ow[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 899.150 53.400 899.450 54.400 ;
    END
  END um_ow[276]
  PIN um_ow[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 895.470 53.400 895.770 54.400 ;
    END
  END um_ow[277]
  PIN um_ow[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 891.790 53.400 892.090 54.400 ;
    END
  END um_ow[278]
  PIN um_ow[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 888.110 53.400 888.410 54.400 ;
    END
  END um_ow[279]
  PIN um_ow[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 53.400 81.570 54.400 ;
    END
  END um_ow[27]
  PIN um_ow[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 884.430 53.400 884.730 54.400 ;
    END
  END um_ow[280]
  PIN um_ow[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 880.750 53.400 881.050 54.400 ;
    END
  END um_ow[281]
  PIN um_ow[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 877.070 53.400 877.370 54.400 ;
    END
  END um_ow[282]
  PIN um_ow[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 873.390 53.400 873.690 54.400 ;
    END
  END um_ow[283]
  PIN um_ow[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 869.710 53.400 870.010 54.400 ;
    END
  END um_ow[284]
  PIN um_ow[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 866.030 53.400 866.330 54.400 ;
    END
  END um_ow[285]
  PIN um_ow[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 862.350 53.400 862.650 54.400 ;
    END
  END um_ow[286]
  PIN um_ow[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 858.670 53.400 858.970 54.400 ;
    END
  END um_ow[287]
  PIN um_ow[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1113.510 0.000 1113.810 1.000 ;
    END
  END um_ow[288]
  PIN um_ow[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1109.830 0.000 1110.130 1.000 ;
    END
  END um_ow[289]
  PIN um_ow[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 53.400 77.890 54.400 ;
    END
  END um_ow[28]
  PIN um_ow[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1106.150 0.000 1106.450 1.000 ;
    END
  END um_ow[290]
  PIN um_ow[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1102.470 0.000 1102.770 1.000 ;
    END
  END um_ow[291]
  PIN um_ow[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1098.790 0.000 1099.090 1.000 ;
    END
  END um_ow[292]
  PIN um_ow[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1095.110 0.000 1095.410 1.000 ;
    END
  END um_ow[293]
  PIN um_ow[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1091.430 0.000 1091.730 1.000 ;
    END
  END um_ow[294]
  PIN um_ow[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1087.750 0.000 1088.050 1.000 ;
    END
  END um_ow[295]
  PIN um_ow[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1084.070 0.000 1084.370 1.000 ;
    END
  END um_ow[296]
  PIN um_ow[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1080.390 0.000 1080.690 1.000 ;
    END
  END um_ow[297]
  PIN um_ow[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1076.710 0.000 1077.010 1.000 ;
    END
  END um_ow[298]
  PIN um_ow[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1073.030 0.000 1073.330 1.000 ;
    END
  END um_ow[299]
  PIN um_ow[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 73.910 53.400 74.210 54.400 ;
    END
  END um_ow[29]
  PIN um_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.950 0.000 85.250 1.000 ;
    END
  END um_ow[2]
  PIN um_ow[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1069.350 0.000 1069.650 1.000 ;
    END
  END um_ow[300]
  PIN um_ow[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1065.670 0.000 1065.970 1.000 ;
    END
  END um_ow[301]
  PIN um_ow[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1061.990 0.000 1062.290 1.000 ;
    END
  END um_ow[302]
  PIN um_ow[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1058.310 0.000 1058.610 1.000 ;
    END
  END um_ow[303]
  PIN um_ow[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1054.630 0.000 1054.930 1.000 ;
    END
  END um_ow[304]
  PIN um_ow[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1050.950 0.000 1051.250 1.000 ;
    END
  END um_ow[305]
  PIN um_ow[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1047.270 0.000 1047.570 1.000 ;
    END
  END um_ow[306]
  PIN um_ow[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1043.590 0.000 1043.890 1.000 ;
    END
  END um_ow[307]
  PIN um_ow[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1039.910 0.000 1040.210 1.000 ;
    END
  END um_ow[308]
  PIN um_ow[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1036.230 0.000 1036.530 1.000 ;
    END
  END um_ow[309]
  PIN um_ow[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 53.400 70.530 54.400 ;
    END
  END um_ow[30]
  PIN um_ow[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1032.550 0.000 1032.850 1.000 ;
    END
  END um_ow[310]
  PIN um_ow[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1028.870 0.000 1029.170 1.000 ;
    END
  END um_ow[311]
  PIN um_ow[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1113.510 53.400 1113.810 54.400 ;
    END
  END um_ow[312]
  PIN um_ow[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1109.830 53.400 1110.130 54.400 ;
    END
  END um_ow[313]
  PIN um_ow[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1106.150 53.400 1106.450 54.400 ;
    END
  END um_ow[314]
  PIN um_ow[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1102.470 53.400 1102.770 54.400 ;
    END
  END um_ow[315]
  PIN um_ow[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1098.790 53.400 1099.090 54.400 ;
    END
  END um_ow[316]
  PIN um_ow[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1095.110 53.400 1095.410 54.400 ;
    END
  END um_ow[317]
  PIN um_ow[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1091.430 53.400 1091.730 54.400 ;
    END
  END um_ow[318]
  PIN um_ow[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1087.750 53.400 1088.050 54.400 ;
    END
  END um_ow[319]
  PIN um_ow[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 53.400 66.850 54.400 ;
    END
  END um_ow[31]
  PIN um_ow[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1084.070 53.400 1084.370 54.400 ;
    END
  END um_ow[320]
  PIN um_ow[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1080.390 53.400 1080.690 54.400 ;
    END
  END um_ow[321]
  PIN um_ow[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1076.710 53.400 1077.010 54.400 ;
    END
  END um_ow[322]
  PIN um_ow[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1073.030 53.400 1073.330 54.400 ;
    END
  END um_ow[323]
  PIN um_ow[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1069.350 53.400 1069.650 54.400 ;
    END
  END um_ow[324]
  PIN um_ow[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1065.670 53.400 1065.970 54.400 ;
    END
  END um_ow[325]
  PIN um_ow[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1061.990 53.400 1062.290 54.400 ;
    END
  END um_ow[326]
  PIN um_ow[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1058.310 53.400 1058.610 54.400 ;
    END
  END um_ow[327]
  PIN um_ow[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1054.630 53.400 1054.930 54.400 ;
    END
  END um_ow[328]
  PIN um_ow[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1050.950 53.400 1051.250 54.400 ;
    END
  END um_ow[329]
  PIN um_ow[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 53.400 63.170 54.400 ;
    END
  END um_ow[32]
  PIN um_ow[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1047.270 53.400 1047.570 54.400 ;
    END
  END um_ow[330]
  PIN um_ow[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1043.590 53.400 1043.890 54.400 ;
    END
  END um_ow[331]
  PIN um_ow[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1039.910 53.400 1040.210 54.400 ;
    END
  END um_ow[332]
  PIN um_ow[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1036.230 53.400 1036.530 54.400 ;
    END
  END um_ow[333]
  PIN um_ow[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1032.550 53.400 1032.850 54.400 ;
    END
  END um_ow[334]
  PIN um_ow[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1028.870 53.400 1029.170 54.400 ;
    END
  END um_ow[335]
  PIN um_ow[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1283.710 0.000 1284.010 1.000 ;
    END
  END um_ow[336]
  PIN um_ow[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1280.030 0.000 1280.330 1.000 ;
    END
  END um_ow[337]
  PIN um_ow[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1276.350 0.000 1276.650 1.000 ;
    END
  END um_ow[338]
  PIN um_ow[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1272.670 0.000 1272.970 1.000 ;
    END
  END um_ow[339]
  PIN um_ow[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 53.400 59.490 54.400 ;
    END
  END um_ow[33]
  PIN um_ow[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1268.990 0.000 1269.290 1.000 ;
    END
  END um_ow[340]
  PIN um_ow[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1265.310 0.000 1265.610 1.000 ;
    END
  END um_ow[341]
  PIN um_ow[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1261.630 0.000 1261.930 1.000 ;
    END
  END um_ow[342]
  PIN um_ow[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1257.950 0.000 1258.250 1.000 ;
    END
  END um_ow[343]
  PIN um_ow[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1254.270 0.000 1254.570 1.000 ;
    END
  END um_ow[344]
  PIN um_ow[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1250.590 0.000 1250.890 1.000 ;
    END
  END um_ow[345]
  PIN um_ow[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1246.910 0.000 1247.210 1.000 ;
    END
  END um_ow[346]
  PIN um_ow[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1243.230 0.000 1243.530 1.000 ;
    END
  END um_ow[347]
  PIN um_ow[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1239.550 0.000 1239.850 1.000 ;
    END
  END um_ow[348]
  PIN um_ow[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1235.870 0.000 1236.170 1.000 ;
    END
  END um_ow[349]
  PIN um_ow[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 53.400 55.810 54.400 ;
    END
  END um_ow[34]
  PIN um_ow[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1232.190 0.000 1232.490 1.000 ;
    END
  END um_ow[350]
  PIN um_ow[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1228.510 0.000 1228.810 1.000 ;
    END
  END um_ow[351]
  PIN um_ow[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1224.830 0.000 1225.130 1.000 ;
    END
  END um_ow[352]
  PIN um_ow[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1221.150 0.000 1221.450 1.000 ;
    END
  END um_ow[353]
  PIN um_ow[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1217.470 0.000 1217.770 1.000 ;
    END
  END um_ow[354]
  PIN um_ow[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1213.790 0.000 1214.090 1.000 ;
    END
  END um_ow[355]
  PIN um_ow[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1210.110 0.000 1210.410 1.000 ;
    END
  END um_ow[356]
  PIN um_ow[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1206.430 0.000 1206.730 1.000 ;
    END
  END um_ow[357]
  PIN um_ow[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1202.750 0.000 1203.050 1.000 ;
    END
  END um_ow[358]
  PIN um_ow[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1199.070 0.000 1199.370 1.000 ;
    END
  END um_ow[359]
  PIN um_ow[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 51.830 53.400 52.130 54.400 ;
    END
  END um_ow[35]
  PIN um_ow[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1283.710 53.400 1284.010 54.400 ;
    END
  END um_ow[360]
  PIN um_ow[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1280.030 53.400 1280.330 54.400 ;
    END
  END um_ow[361]
  PIN um_ow[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1276.350 53.400 1276.650 54.400 ;
    END
  END um_ow[362]
  PIN um_ow[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1272.670 53.400 1272.970 54.400 ;
    END
  END um_ow[363]
  PIN um_ow[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1268.990 53.400 1269.290 54.400 ;
    END
  END um_ow[364]
  PIN um_ow[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1265.310 53.400 1265.610 54.400 ;
    END
  END um_ow[365]
  PIN um_ow[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1261.630 53.400 1261.930 54.400 ;
    END
  END um_ow[366]
  PIN um_ow[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1257.950 53.400 1258.250 54.400 ;
    END
  END um_ow[367]
  PIN um_ow[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1254.270 53.400 1254.570 54.400 ;
    END
  END um_ow[368]
  PIN um_ow[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1250.590 53.400 1250.890 54.400 ;
    END
  END um_ow[369]
  PIN um_ow[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 53.400 48.450 54.400 ;
    END
  END um_ow[36]
  PIN um_ow[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1246.910 53.400 1247.210 54.400 ;
    END
  END um_ow[370]
  PIN um_ow[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1243.230 53.400 1243.530 54.400 ;
    END
  END um_ow[371]
  PIN um_ow[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1239.550 53.400 1239.850 54.400 ;
    END
  END um_ow[372]
  PIN um_ow[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1235.870 53.400 1236.170 54.400 ;
    END
  END um_ow[373]
  PIN um_ow[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1232.190 53.400 1232.490 54.400 ;
    END
  END um_ow[374]
  PIN um_ow[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1228.510 53.400 1228.810 54.400 ;
    END
  END um_ow[375]
  PIN um_ow[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1224.830 53.400 1225.130 54.400 ;
    END
  END um_ow[376]
  PIN um_ow[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1221.150 53.400 1221.450 54.400 ;
    END
  END um_ow[377]
  PIN um_ow[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1217.470 53.400 1217.770 54.400 ;
    END
  END um_ow[378]
  PIN um_ow[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 1213.790 53.400 1214.090 54.400 ;
    END
  END um_ow[379]
  PIN um_ow[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 53.400 44.770 54.400 ;
    END
  END um_ow[37]
  PIN um_ow[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1210.110 53.400 1210.410 54.400 ;
    END
  END um_ow[380]
  PIN um_ow[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1206.430 53.400 1206.730 54.400 ;
    END
  END um_ow[381]
  PIN um_ow[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1202.750 53.400 1203.050 54.400 ;
    END
  END um_ow[382]
  PIN um_ow[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1199.070 53.400 1199.370 54.400 ;
    END
  END um_ow[383]
  PIN um_ow[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 40.790 53.400 41.090 54.400 ;
    END
  END um_ow[38]
  PIN um_ow[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 37.110 53.400 37.410 54.400 ;
    END
  END um_ow[39]
  PIN um_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 81.270 0.000 81.570 1.000 ;
    END
  END um_ow[3]
  PIN um_ow[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 33.430 53.400 33.730 54.400 ;
    END
  END um_ow[40]
  PIN um_ow[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 29.750 53.400 30.050 54.400 ;
    END
  END um_ow[41]
  PIN um_ow[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 53.400 26.370 54.400 ;
    END
  END um_ow[42]
  PIN um_ow[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 22.390 53.400 22.690 54.400 ;
    END
  END um_ow[43]
  PIN um_ow[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 18.710 53.400 19.010 54.400 ;
    END
  END um_ow[44]
  PIN um_ow[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 15.030 53.400 15.330 54.400 ;
    END
  END um_ow[45]
  PIN um_ow[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 11.350 53.400 11.650 54.400 ;
    END
  END um_ow[46]
  PIN um_ow[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 7.670 53.400 7.970 54.400 ;
    END
  END um_ow[47]
  PIN um_ow[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 262.510 0.000 262.810 1.000 ;
    END
  END um_ow[48]
  PIN um_ow[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 258.830 0.000 259.130 1.000 ;
    END
  END um_ow[49]
  PIN um_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 77.590 0.000 77.890 1.000 ;
    END
  END um_ow[4]
  PIN um_ow[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 255.150 0.000 255.450 1.000 ;
    END
  END um_ow[50]
  PIN um_ow[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 251.470 0.000 251.770 1.000 ;
    END
  END um_ow[51]
  PIN um_ow[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 247.790 0.000 248.090 1.000 ;
    END
  END um_ow[52]
  PIN um_ow[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 244.110 0.000 244.410 1.000 ;
    END
  END um_ow[53]
  PIN um_ow[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 240.430 0.000 240.730 1.000 ;
    END
  END um_ow[54]
  PIN um_ow[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 236.750 0.000 237.050 1.000 ;
    END
  END um_ow[55]
  PIN um_ow[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 233.070 0.000 233.370 1.000 ;
    END
  END um_ow[56]
  PIN um_ow[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 229.390 0.000 229.690 1.000 ;
    END
  END um_ow[57]
  PIN um_ow[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 225.710 0.000 226.010 1.000 ;
    END
  END um_ow[58]
  PIN um_ow[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 222.030 0.000 222.330 1.000 ;
    END
  END um_ow[59]
  PIN um_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 73.910 0.000 74.210 1.000 ;
    END
  END um_ow[5]
  PIN um_ow[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 218.350 0.000 218.650 1.000 ;
    END
  END um_ow[60]
  PIN um_ow[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 214.670 0.000 214.970 1.000 ;
    END
  END um_ow[61]
  PIN um_ow[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 210.990 0.000 211.290 1.000 ;
    END
  END um_ow[62]
  PIN um_ow[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 207.310 0.000 207.610 1.000 ;
    END
  END um_ow[63]
  PIN um_ow[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 203.630 0.000 203.930 1.000 ;
    END
  END um_ow[64]
  PIN um_ow[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 199.950 0.000 200.250 1.000 ;
    END
  END um_ow[65]
  PIN um_ow[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 196.270 0.000 196.570 1.000 ;
    END
  END um_ow[66]
  PIN um_ow[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 192.590 0.000 192.890 1.000 ;
    END
  END um_ow[67]
  PIN um_ow[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 188.910 0.000 189.210 1.000 ;
    END
  END um_ow[68]
  PIN um_ow[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 185.230 0.000 185.530 1.000 ;
    END
  END um_ow[69]
  PIN um_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 70.230 0.000 70.530 1.000 ;
    END
  END um_ow[6]
  PIN um_ow[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 181.550 0.000 181.850 1.000 ;
    END
  END um_ow[70]
  PIN um_ow[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 177.870 0.000 178.170 1.000 ;
    END
  END um_ow[71]
  PIN um_ow[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 262.510 53.400 262.810 54.400 ;
    END
  END um_ow[72]
  PIN um_ow[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 258.830 53.400 259.130 54.400 ;
    END
  END um_ow[73]
  PIN um_ow[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 255.150 53.400 255.450 54.400 ;
    END
  END um_ow[74]
  PIN um_ow[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 251.470 53.400 251.770 54.400 ;
    END
  END um_ow[75]
  PIN um_ow[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 247.790 53.400 248.090 54.400 ;
    END
  END um_ow[76]
  PIN um_ow[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 244.110 53.400 244.410 54.400 ;
    END
  END um_ow[77]
  PIN um_ow[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 240.430 53.400 240.730 54.400 ;
    END
  END um_ow[78]
  PIN um_ow[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 236.750 53.400 237.050 54.400 ;
    END
  END um_ow[79]
  PIN um_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 66.550 0.000 66.850 1.000 ;
    END
  END um_ow[7]
  PIN um_ow[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 233.070 53.400 233.370 54.400 ;
    END
  END um_ow[80]
  PIN um_ow[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 229.390 53.400 229.690 54.400 ;
    END
  END um_ow[81]
  PIN um_ow[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 225.710 53.400 226.010 54.400 ;
    END
  END um_ow[82]
  PIN um_ow[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 222.030 53.400 222.330 54.400 ;
    END
  END um_ow[83]
  PIN um_ow[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 218.350 53.400 218.650 54.400 ;
    END
  END um_ow[84]
  PIN um_ow[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 214.670 53.400 214.970 54.400 ;
    END
  END um_ow[85]
  PIN um_ow[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 210.990 53.400 211.290 54.400 ;
    END
  END um_ow[86]
  PIN um_ow[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 207.310 53.400 207.610 54.400 ;
    END
  END um_ow[87]
  PIN um_ow[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 203.630 53.400 203.930 54.400 ;
    END
  END um_ow[88]
  PIN um_ow[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 199.950 53.400 200.250 54.400 ;
    END
  END um_ow[89]
  PIN um_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 0.000 63.170 1.000 ;
    END
  END um_ow[8]
  PIN um_ow[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 196.270 53.400 196.570 54.400 ;
    END
  END um_ow[90]
  PIN um_ow[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 192.590 53.400 192.890 54.400 ;
    END
  END um_ow[91]
  PIN um_ow[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 188.910 53.400 189.210 54.400 ;
    END
  END um_ow[92]
  PIN um_ow[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 185.230 53.400 185.530 54.400 ;
    END
  END um_ow[93]
  PIN um_ow[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 181.550 53.400 181.850 54.400 ;
    END
  END um_ow[94]
  PIN um_ow[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 177.870 53.400 178.170 54.400 ;
    END
  END um_ow[95]
  PIN um_ow[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 432.710 0.000 433.010 1.000 ;
    END
  END um_ow[96]
  PIN um_ow[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 429.030 0.000 429.330 1.000 ;
    END
  END um_ow[97]
  PIN um_ow[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 425.350 0.000 425.650 1.000 ;
    END
  END um_ow[98]
  PIN um_ow[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 421.670 0.000 421.970 1.000 ;
    END
  END um_ow[99]
  PIN um_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 59.190 0.000 59.490 1.000 ;
    END
  END um_ow[9]
  OBS
      LAYER nwell ;
        RECT 2.570 47.545 1356.270 50.375 ;
        RECT 2.570 42.105 1356.270 44.935 ;
        RECT 2.570 36.665 1356.270 39.495 ;
        RECT 2.570 31.225 1356.270 34.055 ;
        RECT 2.570 25.785 1356.270 28.615 ;
        RECT 2.570 20.345 1356.270 23.175 ;
        RECT 2.570 14.905 1356.270 17.735 ;
        RECT 2.570 9.465 1356.270 12.295 ;
        RECT 2.570 4.025 1356.270 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 1356.080 51.765 ;
      LAYER met1 ;
        RECT 2.760 0.040 1356.080 54.360 ;
      LAYER met2 ;
        RECT 4.230 0.010 1355.060 54.390 ;
      LAYER met3 ;
        RECT 3.750 48.490 1357.840 52.865 ;
        RECT 3.750 4.550 1357.440 48.490 ;
        RECT 3.750 0.175 1357.840 4.550 ;
      LAYER met4 ;
        RECT 4.690 53.000 7.270 54.050 ;
        RECT 8.370 53.000 10.950 54.050 ;
        RECT 12.050 53.000 14.630 54.050 ;
        RECT 15.730 53.000 18.310 54.050 ;
        RECT 19.410 53.000 21.990 54.050 ;
        RECT 23.090 53.000 25.670 54.050 ;
        RECT 26.770 53.000 29.350 54.050 ;
        RECT 30.450 53.000 33.030 54.050 ;
        RECT 34.130 53.000 36.710 54.050 ;
        RECT 37.810 53.000 40.390 54.050 ;
        RECT 41.490 53.000 44.070 54.050 ;
        RECT 45.170 53.000 47.750 54.050 ;
        RECT 48.850 53.000 51.430 54.050 ;
        RECT 52.530 53.000 55.110 54.050 ;
        RECT 56.210 53.000 58.790 54.050 ;
        RECT 59.890 53.000 62.470 54.050 ;
        RECT 63.570 53.000 66.150 54.050 ;
        RECT 67.250 53.000 69.830 54.050 ;
        RECT 70.930 53.000 73.510 54.050 ;
        RECT 74.610 53.000 77.190 54.050 ;
        RECT 78.290 53.000 80.870 54.050 ;
        RECT 81.970 53.000 84.550 54.050 ;
        RECT 85.650 53.000 88.230 54.050 ;
        RECT 89.330 53.000 91.910 54.050 ;
        RECT 93.010 53.000 95.590 54.050 ;
        RECT 96.690 53.000 99.270 54.050 ;
        RECT 100.370 53.000 102.950 54.050 ;
        RECT 104.050 53.000 106.630 54.050 ;
        RECT 107.730 53.000 110.310 54.050 ;
        RECT 111.410 53.000 113.990 54.050 ;
        RECT 115.090 53.000 117.670 54.050 ;
        RECT 118.770 53.000 121.350 54.050 ;
        RECT 122.450 53.000 125.030 54.050 ;
        RECT 126.130 53.000 128.710 54.050 ;
        RECT 129.810 53.000 132.390 54.050 ;
        RECT 133.490 53.000 136.070 54.050 ;
        RECT 137.170 53.000 139.750 54.050 ;
        RECT 140.850 53.000 143.430 54.050 ;
        RECT 144.530 53.000 147.110 54.050 ;
        RECT 148.210 53.000 150.790 54.050 ;
        RECT 151.890 53.000 154.470 54.050 ;
        RECT 155.570 53.000 158.150 54.050 ;
        RECT 159.250 53.000 161.830 54.050 ;
        RECT 162.930 53.000 173.790 54.050 ;
        RECT 174.890 53.000 177.470 54.050 ;
        RECT 178.570 53.000 181.150 54.050 ;
        RECT 182.250 53.000 184.830 54.050 ;
        RECT 185.930 53.000 188.510 54.050 ;
        RECT 189.610 53.000 192.190 54.050 ;
        RECT 193.290 53.000 195.870 54.050 ;
        RECT 196.970 53.000 199.550 54.050 ;
        RECT 200.650 53.000 203.230 54.050 ;
        RECT 204.330 53.000 206.910 54.050 ;
        RECT 208.010 53.000 210.590 54.050 ;
        RECT 211.690 53.000 214.270 54.050 ;
        RECT 215.370 53.000 217.950 54.050 ;
        RECT 219.050 53.000 221.630 54.050 ;
        RECT 222.730 53.000 225.310 54.050 ;
        RECT 226.410 53.000 228.990 54.050 ;
        RECT 230.090 53.000 232.670 54.050 ;
        RECT 233.770 53.000 236.350 54.050 ;
        RECT 237.450 53.000 240.030 54.050 ;
        RECT 241.130 53.000 243.710 54.050 ;
        RECT 244.810 53.000 247.390 54.050 ;
        RECT 248.490 53.000 251.070 54.050 ;
        RECT 252.170 53.000 254.750 54.050 ;
        RECT 255.850 53.000 258.430 54.050 ;
        RECT 259.530 53.000 262.110 54.050 ;
        RECT 263.210 53.000 265.790 54.050 ;
        RECT 266.890 53.000 269.470 54.050 ;
        RECT 270.570 53.000 273.150 54.050 ;
        RECT 274.250 53.000 276.830 54.050 ;
        RECT 277.930 53.000 280.510 54.050 ;
        RECT 281.610 53.000 284.190 54.050 ;
        RECT 285.290 53.000 287.870 54.050 ;
        RECT 288.970 53.000 291.550 54.050 ;
        RECT 292.650 53.000 295.230 54.050 ;
        RECT 296.330 53.000 298.910 54.050 ;
        RECT 300.010 53.000 302.590 54.050 ;
        RECT 303.690 53.000 306.270 54.050 ;
        RECT 307.370 53.000 309.950 54.050 ;
        RECT 311.050 53.000 313.630 54.050 ;
        RECT 314.730 53.000 317.310 54.050 ;
        RECT 318.410 53.000 320.990 54.050 ;
        RECT 322.090 53.000 324.670 54.050 ;
        RECT 325.770 53.000 328.350 54.050 ;
        RECT 329.450 53.000 332.030 54.050 ;
        RECT 333.130 53.000 343.990 54.050 ;
        RECT 345.090 53.000 347.670 54.050 ;
        RECT 348.770 53.000 351.350 54.050 ;
        RECT 352.450 53.000 355.030 54.050 ;
        RECT 356.130 53.000 358.710 54.050 ;
        RECT 359.810 53.000 362.390 54.050 ;
        RECT 363.490 53.000 366.070 54.050 ;
        RECT 367.170 53.000 369.750 54.050 ;
        RECT 370.850 53.000 373.430 54.050 ;
        RECT 374.530 53.000 377.110 54.050 ;
        RECT 378.210 53.000 380.790 54.050 ;
        RECT 381.890 53.000 384.470 54.050 ;
        RECT 385.570 53.000 388.150 54.050 ;
        RECT 389.250 53.000 391.830 54.050 ;
        RECT 392.930 53.000 395.510 54.050 ;
        RECT 396.610 53.000 399.190 54.050 ;
        RECT 400.290 53.000 402.870 54.050 ;
        RECT 403.970 53.000 406.550 54.050 ;
        RECT 407.650 53.000 410.230 54.050 ;
        RECT 411.330 53.000 413.910 54.050 ;
        RECT 415.010 53.000 417.590 54.050 ;
        RECT 418.690 53.000 421.270 54.050 ;
        RECT 422.370 53.000 424.950 54.050 ;
        RECT 426.050 53.000 428.630 54.050 ;
        RECT 429.730 53.000 432.310 54.050 ;
        RECT 433.410 53.000 435.990 54.050 ;
        RECT 437.090 53.000 439.670 54.050 ;
        RECT 440.770 53.000 443.350 54.050 ;
        RECT 444.450 53.000 447.030 54.050 ;
        RECT 448.130 53.000 450.710 54.050 ;
        RECT 451.810 53.000 454.390 54.050 ;
        RECT 455.490 53.000 458.070 54.050 ;
        RECT 459.170 53.000 461.750 54.050 ;
        RECT 462.850 53.000 465.430 54.050 ;
        RECT 466.530 53.000 469.110 54.050 ;
        RECT 470.210 53.000 472.790 54.050 ;
        RECT 473.890 53.000 476.470 54.050 ;
        RECT 477.570 53.000 480.150 54.050 ;
        RECT 481.250 53.000 483.830 54.050 ;
        RECT 484.930 53.000 487.510 54.050 ;
        RECT 488.610 53.000 491.190 54.050 ;
        RECT 492.290 53.000 494.870 54.050 ;
        RECT 495.970 53.000 498.550 54.050 ;
        RECT 499.650 53.000 502.230 54.050 ;
        RECT 503.330 53.000 514.190 54.050 ;
        RECT 515.290 53.000 517.870 54.050 ;
        RECT 518.970 53.000 521.550 54.050 ;
        RECT 522.650 53.000 525.230 54.050 ;
        RECT 526.330 53.000 528.910 54.050 ;
        RECT 530.010 53.000 532.590 54.050 ;
        RECT 533.690 53.000 536.270 54.050 ;
        RECT 537.370 53.000 539.950 54.050 ;
        RECT 541.050 53.000 543.630 54.050 ;
        RECT 544.730 53.000 547.310 54.050 ;
        RECT 548.410 53.000 550.990 54.050 ;
        RECT 552.090 53.000 554.670 54.050 ;
        RECT 555.770 53.000 558.350 54.050 ;
        RECT 559.450 53.000 562.030 54.050 ;
        RECT 563.130 53.000 565.710 54.050 ;
        RECT 566.810 53.000 569.390 54.050 ;
        RECT 570.490 53.000 573.070 54.050 ;
        RECT 574.170 53.000 576.750 54.050 ;
        RECT 577.850 53.000 580.430 54.050 ;
        RECT 581.530 53.000 584.110 54.050 ;
        RECT 585.210 53.000 587.790 54.050 ;
        RECT 588.890 53.000 591.470 54.050 ;
        RECT 592.570 53.000 595.150 54.050 ;
        RECT 596.250 53.000 598.830 54.050 ;
        RECT 599.930 53.000 602.510 54.050 ;
        RECT 603.610 53.000 606.190 54.050 ;
        RECT 607.290 53.000 609.870 54.050 ;
        RECT 610.970 53.000 613.550 54.050 ;
        RECT 614.650 53.000 617.230 54.050 ;
        RECT 618.330 53.000 620.910 54.050 ;
        RECT 622.010 53.000 624.590 54.050 ;
        RECT 625.690 53.000 628.270 54.050 ;
        RECT 629.370 53.000 631.950 54.050 ;
        RECT 633.050 53.000 635.630 54.050 ;
        RECT 636.730 53.000 639.310 54.050 ;
        RECT 640.410 53.000 642.990 54.050 ;
        RECT 644.090 53.000 646.670 54.050 ;
        RECT 647.770 53.000 650.350 54.050 ;
        RECT 651.450 53.000 654.030 54.050 ;
        RECT 655.130 53.000 657.710 54.050 ;
        RECT 658.810 53.000 661.390 54.050 ;
        RECT 662.490 53.000 665.070 54.050 ;
        RECT 666.170 53.000 668.750 54.050 ;
        RECT 669.850 53.000 672.430 54.050 ;
        RECT 673.530 53.000 684.390 54.050 ;
        RECT 685.490 53.000 688.070 54.050 ;
        RECT 689.170 53.000 691.750 54.050 ;
        RECT 692.850 53.000 695.430 54.050 ;
        RECT 696.530 53.000 699.110 54.050 ;
        RECT 700.210 53.000 702.790 54.050 ;
        RECT 703.890 53.000 706.470 54.050 ;
        RECT 707.570 53.000 710.150 54.050 ;
        RECT 711.250 53.000 713.830 54.050 ;
        RECT 714.930 53.000 717.510 54.050 ;
        RECT 718.610 53.000 721.190 54.050 ;
        RECT 722.290 53.000 724.870 54.050 ;
        RECT 725.970 53.000 728.550 54.050 ;
        RECT 729.650 53.000 732.230 54.050 ;
        RECT 733.330 53.000 735.910 54.050 ;
        RECT 737.010 53.000 739.590 54.050 ;
        RECT 740.690 53.000 743.270 54.050 ;
        RECT 744.370 53.000 746.950 54.050 ;
        RECT 748.050 53.000 750.630 54.050 ;
        RECT 751.730 53.000 754.310 54.050 ;
        RECT 755.410 53.000 757.990 54.050 ;
        RECT 759.090 53.000 761.670 54.050 ;
        RECT 762.770 53.000 765.350 54.050 ;
        RECT 766.450 53.000 769.030 54.050 ;
        RECT 770.130 53.000 772.710 54.050 ;
        RECT 773.810 53.000 776.390 54.050 ;
        RECT 777.490 53.000 780.070 54.050 ;
        RECT 781.170 53.000 783.750 54.050 ;
        RECT 784.850 53.000 787.430 54.050 ;
        RECT 788.530 53.000 791.110 54.050 ;
        RECT 792.210 53.000 794.790 54.050 ;
        RECT 795.890 53.000 798.470 54.050 ;
        RECT 799.570 53.000 802.150 54.050 ;
        RECT 803.250 53.000 805.830 54.050 ;
        RECT 806.930 53.000 809.510 54.050 ;
        RECT 810.610 53.000 813.190 54.050 ;
        RECT 814.290 53.000 816.870 54.050 ;
        RECT 817.970 53.000 820.550 54.050 ;
        RECT 821.650 53.000 824.230 54.050 ;
        RECT 825.330 53.000 827.910 54.050 ;
        RECT 829.010 53.000 831.590 54.050 ;
        RECT 832.690 53.000 835.270 54.050 ;
        RECT 836.370 53.000 838.950 54.050 ;
        RECT 840.050 53.000 842.630 54.050 ;
        RECT 843.730 53.000 854.590 54.050 ;
        RECT 855.690 53.000 858.270 54.050 ;
        RECT 859.370 53.000 861.950 54.050 ;
        RECT 863.050 53.000 865.630 54.050 ;
        RECT 866.730 53.000 869.310 54.050 ;
        RECT 870.410 53.000 872.990 54.050 ;
        RECT 874.090 53.000 876.670 54.050 ;
        RECT 877.770 53.000 880.350 54.050 ;
        RECT 881.450 53.000 884.030 54.050 ;
        RECT 885.130 53.000 887.710 54.050 ;
        RECT 888.810 53.000 891.390 54.050 ;
        RECT 892.490 53.000 895.070 54.050 ;
        RECT 896.170 53.000 898.750 54.050 ;
        RECT 899.850 53.000 902.430 54.050 ;
        RECT 903.530 53.000 906.110 54.050 ;
        RECT 907.210 53.000 909.790 54.050 ;
        RECT 910.890 53.000 913.470 54.050 ;
        RECT 914.570 53.000 917.150 54.050 ;
        RECT 918.250 53.000 920.830 54.050 ;
        RECT 921.930 53.000 924.510 54.050 ;
        RECT 925.610 53.000 928.190 54.050 ;
        RECT 929.290 53.000 931.870 54.050 ;
        RECT 932.970 53.000 935.550 54.050 ;
        RECT 936.650 53.000 939.230 54.050 ;
        RECT 940.330 53.000 942.910 54.050 ;
        RECT 944.010 53.000 946.590 54.050 ;
        RECT 947.690 53.000 950.270 54.050 ;
        RECT 951.370 53.000 953.950 54.050 ;
        RECT 955.050 53.000 957.630 54.050 ;
        RECT 958.730 53.000 961.310 54.050 ;
        RECT 962.410 53.000 964.990 54.050 ;
        RECT 966.090 53.000 968.670 54.050 ;
        RECT 969.770 53.000 972.350 54.050 ;
        RECT 973.450 53.000 976.030 54.050 ;
        RECT 977.130 53.000 979.710 54.050 ;
        RECT 980.810 53.000 983.390 54.050 ;
        RECT 984.490 53.000 987.070 54.050 ;
        RECT 988.170 53.000 990.750 54.050 ;
        RECT 991.850 53.000 994.430 54.050 ;
        RECT 995.530 53.000 998.110 54.050 ;
        RECT 999.210 53.000 1001.790 54.050 ;
        RECT 1002.890 53.000 1005.470 54.050 ;
        RECT 1006.570 53.000 1009.150 54.050 ;
        RECT 1010.250 53.000 1012.830 54.050 ;
        RECT 1013.930 53.000 1024.790 54.050 ;
        RECT 1025.890 53.000 1028.470 54.050 ;
        RECT 1029.570 53.000 1032.150 54.050 ;
        RECT 1033.250 53.000 1035.830 54.050 ;
        RECT 1036.930 53.000 1039.510 54.050 ;
        RECT 1040.610 53.000 1043.190 54.050 ;
        RECT 1044.290 53.000 1046.870 54.050 ;
        RECT 1047.970 53.000 1050.550 54.050 ;
        RECT 1051.650 53.000 1054.230 54.050 ;
        RECT 1055.330 53.000 1057.910 54.050 ;
        RECT 1059.010 53.000 1061.590 54.050 ;
        RECT 1062.690 53.000 1065.270 54.050 ;
        RECT 1066.370 53.000 1068.950 54.050 ;
        RECT 1070.050 53.000 1072.630 54.050 ;
        RECT 1073.730 53.000 1076.310 54.050 ;
        RECT 1077.410 53.000 1079.990 54.050 ;
        RECT 1081.090 53.000 1083.670 54.050 ;
        RECT 1084.770 53.000 1087.350 54.050 ;
        RECT 1088.450 53.000 1091.030 54.050 ;
        RECT 1092.130 53.000 1094.710 54.050 ;
        RECT 1095.810 53.000 1098.390 54.050 ;
        RECT 1099.490 53.000 1102.070 54.050 ;
        RECT 1103.170 53.000 1105.750 54.050 ;
        RECT 1106.850 53.000 1109.430 54.050 ;
        RECT 1110.530 53.000 1113.110 54.050 ;
        RECT 1114.210 53.000 1116.790 54.050 ;
        RECT 1117.890 53.000 1120.470 54.050 ;
        RECT 1121.570 53.000 1124.150 54.050 ;
        RECT 1125.250 53.000 1127.830 54.050 ;
        RECT 1128.930 53.000 1131.510 54.050 ;
        RECT 1132.610 53.000 1135.190 54.050 ;
        RECT 1136.290 53.000 1138.870 54.050 ;
        RECT 1139.970 53.000 1142.550 54.050 ;
        RECT 1143.650 53.000 1146.230 54.050 ;
        RECT 1147.330 53.000 1149.910 54.050 ;
        RECT 1151.010 53.000 1153.590 54.050 ;
        RECT 1154.690 53.000 1157.270 54.050 ;
        RECT 1158.370 53.000 1160.950 54.050 ;
        RECT 1162.050 53.000 1164.630 54.050 ;
        RECT 1165.730 53.000 1168.310 54.050 ;
        RECT 1169.410 53.000 1171.990 54.050 ;
        RECT 1173.090 53.000 1175.670 54.050 ;
        RECT 1176.770 53.000 1179.350 54.050 ;
        RECT 1180.450 53.000 1183.030 54.050 ;
        RECT 1184.130 53.000 1194.990 54.050 ;
        RECT 1196.090 53.000 1198.670 54.050 ;
        RECT 1199.770 53.000 1202.350 54.050 ;
        RECT 1203.450 53.000 1206.030 54.050 ;
        RECT 1207.130 53.000 1209.710 54.050 ;
        RECT 1210.810 53.000 1213.390 54.050 ;
        RECT 1214.490 53.000 1217.070 54.050 ;
        RECT 1218.170 53.000 1220.750 54.050 ;
        RECT 1221.850 53.000 1224.430 54.050 ;
        RECT 1225.530 53.000 1228.110 54.050 ;
        RECT 1229.210 53.000 1231.790 54.050 ;
        RECT 1232.890 53.000 1235.470 54.050 ;
        RECT 1236.570 53.000 1239.150 54.050 ;
        RECT 1240.250 53.000 1242.830 54.050 ;
        RECT 1243.930 53.000 1246.510 54.050 ;
        RECT 1247.610 53.000 1250.190 54.050 ;
        RECT 1251.290 53.000 1253.870 54.050 ;
        RECT 1254.970 53.000 1257.550 54.050 ;
        RECT 1258.650 53.000 1261.230 54.050 ;
        RECT 1262.330 53.000 1264.910 54.050 ;
        RECT 1266.010 53.000 1268.590 54.050 ;
        RECT 1269.690 53.000 1272.270 54.050 ;
        RECT 1273.370 53.000 1275.950 54.050 ;
        RECT 1277.050 53.000 1279.630 54.050 ;
        RECT 1280.730 53.000 1283.310 54.050 ;
        RECT 1284.410 53.000 1286.990 54.050 ;
        RECT 1288.090 53.000 1290.670 54.050 ;
        RECT 1291.770 53.000 1294.350 54.050 ;
        RECT 1295.450 53.000 1298.030 54.050 ;
        RECT 1299.130 53.000 1301.710 54.050 ;
        RECT 1302.810 53.000 1305.390 54.050 ;
        RECT 1306.490 53.000 1309.070 54.050 ;
        RECT 1310.170 53.000 1312.750 54.050 ;
        RECT 1313.850 53.000 1316.430 54.050 ;
        RECT 1317.530 53.000 1320.110 54.050 ;
        RECT 1321.210 53.000 1323.790 54.050 ;
        RECT 1324.890 53.000 1327.470 54.050 ;
        RECT 1328.570 53.000 1331.150 54.050 ;
        RECT 1332.250 53.000 1334.830 54.050 ;
        RECT 1335.930 53.000 1338.510 54.050 ;
        RECT 1339.610 53.000 1342.190 54.050 ;
        RECT 1343.290 53.000 1345.870 54.050 ;
        RECT 1346.970 53.000 1349.550 54.050 ;
        RECT 1350.650 53.000 1353.230 54.050 ;
        RECT 3.975 52.320 1353.930 53.000 ;
        RECT 3.975 2.080 17.880 52.320 ;
        RECT 20.280 2.080 94.680 52.320 ;
        RECT 97.080 2.080 171.480 52.320 ;
        RECT 173.880 2.080 248.280 52.320 ;
        RECT 250.680 2.080 325.080 52.320 ;
        RECT 327.480 2.080 401.880 52.320 ;
        RECT 404.280 2.080 478.680 52.320 ;
        RECT 481.080 2.080 555.480 52.320 ;
        RECT 557.880 2.080 632.280 52.320 ;
        RECT 634.680 2.080 709.080 52.320 ;
        RECT 711.480 2.080 785.880 52.320 ;
        RECT 788.280 2.080 862.680 52.320 ;
        RECT 865.080 2.080 939.480 52.320 ;
        RECT 941.880 2.080 1016.280 52.320 ;
        RECT 1018.680 2.080 1093.080 52.320 ;
        RECT 1095.480 2.080 1169.880 52.320 ;
        RECT 1172.280 2.080 1246.680 52.320 ;
        RECT 1249.080 2.080 1323.480 52.320 ;
        RECT 1325.880 2.080 1353.930 52.320 ;
        RECT 3.975 1.400 1353.930 2.080 ;
        RECT 4.690 0.350 7.270 1.400 ;
        RECT 8.370 0.350 10.950 1.400 ;
        RECT 12.050 0.350 14.630 1.400 ;
        RECT 15.730 0.350 18.310 1.400 ;
        RECT 19.410 0.350 21.990 1.400 ;
        RECT 23.090 0.350 25.670 1.400 ;
        RECT 26.770 0.350 29.350 1.400 ;
        RECT 30.450 0.350 33.030 1.400 ;
        RECT 34.130 0.350 36.710 1.400 ;
        RECT 37.810 0.350 40.390 1.400 ;
        RECT 41.490 0.350 44.070 1.400 ;
        RECT 45.170 0.350 47.750 1.400 ;
        RECT 48.850 0.350 51.430 1.400 ;
        RECT 52.530 0.350 55.110 1.400 ;
        RECT 56.210 0.350 58.790 1.400 ;
        RECT 59.890 0.350 62.470 1.400 ;
        RECT 63.570 0.350 66.150 1.400 ;
        RECT 67.250 0.350 69.830 1.400 ;
        RECT 70.930 0.350 73.510 1.400 ;
        RECT 74.610 0.350 77.190 1.400 ;
        RECT 78.290 0.350 80.870 1.400 ;
        RECT 81.970 0.350 84.550 1.400 ;
        RECT 85.650 0.350 88.230 1.400 ;
        RECT 89.330 0.350 91.910 1.400 ;
        RECT 93.010 0.350 95.590 1.400 ;
        RECT 96.690 0.350 99.270 1.400 ;
        RECT 100.370 0.350 102.950 1.400 ;
        RECT 104.050 0.350 106.630 1.400 ;
        RECT 107.730 0.350 110.310 1.400 ;
        RECT 111.410 0.350 113.990 1.400 ;
        RECT 115.090 0.350 117.670 1.400 ;
        RECT 118.770 0.350 121.350 1.400 ;
        RECT 122.450 0.350 125.030 1.400 ;
        RECT 126.130 0.350 128.710 1.400 ;
        RECT 129.810 0.350 132.390 1.400 ;
        RECT 133.490 0.350 136.070 1.400 ;
        RECT 137.170 0.350 139.750 1.400 ;
        RECT 140.850 0.350 143.430 1.400 ;
        RECT 144.530 0.350 147.110 1.400 ;
        RECT 148.210 0.350 150.790 1.400 ;
        RECT 151.890 0.350 154.470 1.400 ;
        RECT 155.570 0.350 158.150 1.400 ;
        RECT 159.250 0.350 161.830 1.400 ;
        RECT 162.930 0.350 173.790 1.400 ;
        RECT 174.890 0.350 177.470 1.400 ;
        RECT 178.570 0.350 181.150 1.400 ;
        RECT 182.250 0.350 184.830 1.400 ;
        RECT 185.930 0.350 188.510 1.400 ;
        RECT 189.610 0.350 192.190 1.400 ;
        RECT 193.290 0.350 195.870 1.400 ;
        RECT 196.970 0.350 199.550 1.400 ;
        RECT 200.650 0.350 203.230 1.400 ;
        RECT 204.330 0.350 206.910 1.400 ;
        RECT 208.010 0.350 210.590 1.400 ;
        RECT 211.690 0.350 214.270 1.400 ;
        RECT 215.370 0.350 217.950 1.400 ;
        RECT 219.050 0.350 221.630 1.400 ;
        RECT 222.730 0.350 225.310 1.400 ;
        RECT 226.410 0.350 228.990 1.400 ;
        RECT 230.090 0.350 232.670 1.400 ;
        RECT 233.770 0.350 236.350 1.400 ;
        RECT 237.450 0.350 240.030 1.400 ;
        RECT 241.130 0.350 243.710 1.400 ;
        RECT 244.810 0.350 247.390 1.400 ;
        RECT 248.490 0.350 251.070 1.400 ;
        RECT 252.170 0.350 254.750 1.400 ;
        RECT 255.850 0.350 258.430 1.400 ;
        RECT 259.530 0.350 262.110 1.400 ;
        RECT 263.210 0.350 265.790 1.400 ;
        RECT 266.890 0.350 269.470 1.400 ;
        RECT 270.570 0.350 273.150 1.400 ;
        RECT 274.250 0.350 276.830 1.400 ;
        RECT 277.930 0.350 280.510 1.400 ;
        RECT 281.610 0.350 284.190 1.400 ;
        RECT 285.290 0.350 287.870 1.400 ;
        RECT 288.970 0.350 291.550 1.400 ;
        RECT 292.650 0.350 295.230 1.400 ;
        RECT 296.330 0.350 298.910 1.400 ;
        RECT 300.010 0.350 302.590 1.400 ;
        RECT 303.690 0.350 306.270 1.400 ;
        RECT 307.370 0.350 309.950 1.400 ;
        RECT 311.050 0.350 313.630 1.400 ;
        RECT 314.730 0.350 317.310 1.400 ;
        RECT 318.410 0.350 320.990 1.400 ;
        RECT 322.090 0.350 324.670 1.400 ;
        RECT 325.770 0.350 328.350 1.400 ;
        RECT 329.450 0.350 332.030 1.400 ;
        RECT 333.130 0.350 343.990 1.400 ;
        RECT 345.090 0.350 347.670 1.400 ;
        RECT 348.770 0.350 351.350 1.400 ;
        RECT 352.450 0.350 355.030 1.400 ;
        RECT 356.130 0.350 358.710 1.400 ;
        RECT 359.810 0.350 362.390 1.400 ;
        RECT 363.490 0.350 366.070 1.400 ;
        RECT 367.170 0.350 369.750 1.400 ;
        RECT 370.850 0.350 373.430 1.400 ;
        RECT 374.530 0.350 377.110 1.400 ;
        RECT 378.210 0.350 380.790 1.400 ;
        RECT 381.890 0.350 384.470 1.400 ;
        RECT 385.570 0.350 388.150 1.400 ;
        RECT 389.250 0.350 391.830 1.400 ;
        RECT 392.930 0.350 395.510 1.400 ;
        RECT 396.610 0.350 399.190 1.400 ;
        RECT 400.290 0.350 402.870 1.400 ;
        RECT 403.970 0.350 406.550 1.400 ;
        RECT 407.650 0.350 410.230 1.400 ;
        RECT 411.330 0.350 413.910 1.400 ;
        RECT 415.010 0.350 417.590 1.400 ;
        RECT 418.690 0.350 421.270 1.400 ;
        RECT 422.370 0.350 424.950 1.400 ;
        RECT 426.050 0.350 428.630 1.400 ;
        RECT 429.730 0.350 432.310 1.400 ;
        RECT 433.410 0.350 435.990 1.400 ;
        RECT 437.090 0.350 439.670 1.400 ;
        RECT 440.770 0.350 443.350 1.400 ;
        RECT 444.450 0.350 447.030 1.400 ;
        RECT 448.130 0.350 450.710 1.400 ;
        RECT 451.810 0.350 454.390 1.400 ;
        RECT 455.490 0.350 458.070 1.400 ;
        RECT 459.170 0.350 461.750 1.400 ;
        RECT 462.850 0.350 465.430 1.400 ;
        RECT 466.530 0.350 469.110 1.400 ;
        RECT 470.210 0.350 472.790 1.400 ;
        RECT 473.890 0.350 476.470 1.400 ;
        RECT 477.570 0.350 480.150 1.400 ;
        RECT 481.250 0.350 483.830 1.400 ;
        RECT 484.930 0.350 487.510 1.400 ;
        RECT 488.610 0.350 491.190 1.400 ;
        RECT 492.290 0.350 494.870 1.400 ;
        RECT 495.970 0.350 498.550 1.400 ;
        RECT 499.650 0.350 502.230 1.400 ;
        RECT 503.330 0.350 514.190 1.400 ;
        RECT 515.290 0.350 517.870 1.400 ;
        RECT 518.970 0.350 521.550 1.400 ;
        RECT 522.650 0.350 525.230 1.400 ;
        RECT 526.330 0.350 528.910 1.400 ;
        RECT 530.010 0.350 532.590 1.400 ;
        RECT 533.690 0.350 536.270 1.400 ;
        RECT 537.370 0.350 539.950 1.400 ;
        RECT 541.050 0.350 543.630 1.400 ;
        RECT 544.730 0.350 547.310 1.400 ;
        RECT 548.410 0.350 550.990 1.400 ;
        RECT 552.090 0.350 554.670 1.400 ;
        RECT 555.770 0.350 558.350 1.400 ;
        RECT 559.450 0.350 562.030 1.400 ;
        RECT 563.130 0.350 565.710 1.400 ;
        RECT 566.810 0.350 569.390 1.400 ;
        RECT 570.490 0.350 573.070 1.400 ;
        RECT 574.170 0.350 576.750 1.400 ;
        RECT 577.850 0.350 580.430 1.400 ;
        RECT 581.530 0.350 584.110 1.400 ;
        RECT 585.210 0.350 587.790 1.400 ;
        RECT 588.890 0.350 591.470 1.400 ;
        RECT 592.570 0.350 595.150 1.400 ;
        RECT 596.250 0.350 598.830 1.400 ;
        RECT 599.930 0.350 602.510 1.400 ;
        RECT 603.610 0.350 606.190 1.400 ;
        RECT 607.290 0.350 609.870 1.400 ;
        RECT 610.970 0.350 613.550 1.400 ;
        RECT 614.650 0.350 617.230 1.400 ;
        RECT 618.330 0.350 620.910 1.400 ;
        RECT 622.010 0.350 624.590 1.400 ;
        RECT 625.690 0.350 628.270 1.400 ;
        RECT 629.370 0.350 631.950 1.400 ;
        RECT 633.050 0.350 635.630 1.400 ;
        RECT 636.730 0.350 639.310 1.400 ;
        RECT 640.410 0.350 642.990 1.400 ;
        RECT 644.090 0.350 646.670 1.400 ;
        RECT 647.770 0.350 650.350 1.400 ;
        RECT 651.450 0.350 654.030 1.400 ;
        RECT 655.130 0.350 657.710 1.400 ;
        RECT 658.810 0.350 661.390 1.400 ;
        RECT 662.490 0.350 665.070 1.400 ;
        RECT 666.170 0.350 668.750 1.400 ;
        RECT 669.850 0.350 672.430 1.400 ;
        RECT 673.530 0.350 684.390 1.400 ;
        RECT 685.490 0.350 688.070 1.400 ;
        RECT 689.170 0.350 691.750 1.400 ;
        RECT 692.850 0.350 695.430 1.400 ;
        RECT 696.530 0.350 699.110 1.400 ;
        RECT 700.210 0.350 702.790 1.400 ;
        RECT 703.890 0.350 706.470 1.400 ;
        RECT 707.570 0.350 710.150 1.400 ;
        RECT 711.250 0.350 713.830 1.400 ;
        RECT 714.930 0.350 717.510 1.400 ;
        RECT 718.610 0.350 721.190 1.400 ;
        RECT 722.290 0.350 724.870 1.400 ;
        RECT 725.970 0.350 728.550 1.400 ;
        RECT 729.650 0.350 732.230 1.400 ;
        RECT 733.330 0.350 735.910 1.400 ;
        RECT 737.010 0.350 739.590 1.400 ;
        RECT 740.690 0.350 743.270 1.400 ;
        RECT 744.370 0.350 746.950 1.400 ;
        RECT 748.050 0.350 750.630 1.400 ;
        RECT 751.730 0.350 754.310 1.400 ;
        RECT 755.410 0.350 757.990 1.400 ;
        RECT 759.090 0.350 761.670 1.400 ;
        RECT 762.770 0.350 765.350 1.400 ;
        RECT 766.450 0.350 769.030 1.400 ;
        RECT 770.130 0.350 772.710 1.400 ;
        RECT 773.810 0.350 776.390 1.400 ;
        RECT 777.490 0.350 780.070 1.400 ;
        RECT 781.170 0.350 783.750 1.400 ;
        RECT 784.850 0.350 787.430 1.400 ;
        RECT 788.530 0.350 791.110 1.400 ;
        RECT 792.210 0.350 794.790 1.400 ;
        RECT 795.890 0.350 798.470 1.400 ;
        RECT 799.570 0.350 802.150 1.400 ;
        RECT 803.250 0.350 805.830 1.400 ;
        RECT 806.930 0.350 809.510 1.400 ;
        RECT 810.610 0.350 813.190 1.400 ;
        RECT 814.290 0.350 816.870 1.400 ;
        RECT 817.970 0.350 820.550 1.400 ;
        RECT 821.650 0.350 824.230 1.400 ;
        RECT 825.330 0.350 827.910 1.400 ;
        RECT 829.010 0.350 831.590 1.400 ;
        RECT 832.690 0.350 835.270 1.400 ;
        RECT 836.370 0.350 838.950 1.400 ;
        RECT 840.050 0.350 842.630 1.400 ;
        RECT 843.730 0.350 854.590 1.400 ;
        RECT 855.690 0.350 858.270 1.400 ;
        RECT 859.370 0.350 861.950 1.400 ;
        RECT 863.050 0.350 865.630 1.400 ;
        RECT 866.730 0.350 869.310 1.400 ;
        RECT 870.410 0.350 872.990 1.400 ;
        RECT 874.090 0.350 876.670 1.400 ;
        RECT 877.770 0.350 880.350 1.400 ;
        RECT 881.450 0.350 884.030 1.400 ;
        RECT 885.130 0.350 887.710 1.400 ;
        RECT 888.810 0.350 891.390 1.400 ;
        RECT 892.490 0.350 895.070 1.400 ;
        RECT 896.170 0.350 898.750 1.400 ;
        RECT 899.850 0.350 902.430 1.400 ;
        RECT 903.530 0.350 906.110 1.400 ;
        RECT 907.210 0.350 909.790 1.400 ;
        RECT 910.890 0.350 913.470 1.400 ;
        RECT 914.570 0.350 917.150 1.400 ;
        RECT 918.250 0.350 920.830 1.400 ;
        RECT 921.930 0.350 924.510 1.400 ;
        RECT 925.610 0.350 928.190 1.400 ;
        RECT 929.290 0.350 931.870 1.400 ;
        RECT 932.970 0.350 935.550 1.400 ;
        RECT 936.650 0.350 939.230 1.400 ;
        RECT 940.330 0.350 942.910 1.400 ;
        RECT 944.010 0.350 946.590 1.400 ;
        RECT 947.690 0.350 950.270 1.400 ;
        RECT 951.370 0.350 953.950 1.400 ;
        RECT 955.050 0.350 957.630 1.400 ;
        RECT 958.730 0.350 961.310 1.400 ;
        RECT 962.410 0.350 964.990 1.400 ;
        RECT 966.090 0.350 968.670 1.400 ;
        RECT 969.770 0.350 972.350 1.400 ;
        RECT 973.450 0.350 976.030 1.400 ;
        RECT 977.130 0.350 979.710 1.400 ;
        RECT 980.810 0.350 983.390 1.400 ;
        RECT 984.490 0.350 987.070 1.400 ;
        RECT 988.170 0.350 990.750 1.400 ;
        RECT 991.850 0.350 994.430 1.400 ;
        RECT 995.530 0.350 998.110 1.400 ;
        RECT 999.210 0.350 1001.790 1.400 ;
        RECT 1002.890 0.350 1005.470 1.400 ;
        RECT 1006.570 0.350 1009.150 1.400 ;
        RECT 1010.250 0.350 1012.830 1.400 ;
        RECT 1013.930 0.350 1024.790 1.400 ;
        RECT 1025.890 0.350 1028.470 1.400 ;
        RECT 1029.570 0.350 1032.150 1.400 ;
        RECT 1033.250 0.350 1035.830 1.400 ;
        RECT 1036.930 0.350 1039.510 1.400 ;
        RECT 1040.610 0.350 1043.190 1.400 ;
        RECT 1044.290 0.350 1046.870 1.400 ;
        RECT 1047.970 0.350 1050.550 1.400 ;
        RECT 1051.650 0.350 1054.230 1.400 ;
        RECT 1055.330 0.350 1057.910 1.400 ;
        RECT 1059.010 0.350 1061.590 1.400 ;
        RECT 1062.690 0.350 1065.270 1.400 ;
        RECT 1066.370 0.350 1068.950 1.400 ;
        RECT 1070.050 0.350 1072.630 1.400 ;
        RECT 1073.730 0.350 1076.310 1.400 ;
        RECT 1077.410 0.350 1079.990 1.400 ;
        RECT 1081.090 0.350 1083.670 1.400 ;
        RECT 1084.770 0.350 1087.350 1.400 ;
        RECT 1088.450 0.350 1091.030 1.400 ;
        RECT 1092.130 0.350 1094.710 1.400 ;
        RECT 1095.810 0.350 1098.390 1.400 ;
        RECT 1099.490 0.350 1102.070 1.400 ;
        RECT 1103.170 0.350 1105.750 1.400 ;
        RECT 1106.850 0.350 1109.430 1.400 ;
        RECT 1110.530 0.350 1113.110 1.400 ;
        RECT 1114.210 0.350 1116.790 1.400 ;
        RECT 1117.890 0.350 1120.470 1.400 ;
        RECT 1121.570 0.350 1124.150 1.400 ;
        RECT 1125.250 0.350 1127.830 1.400 ;
        RECT 1128.930 0.350 1131.510 1.400 ;
        RECT 1132.610 0.350 1135.190 1.400 ;
        RECT 1136.290 0.350 1138.870 1.400 ;
        RECT 1139.970 0.350 1142.550 1.400 ;
        RECT 1143.650 0.350 1146.230 1.400 ;
        RECT 1147.330 0.350 1149.910 1.400 ;
        RECT 1151.010 0.350 1153.590 1.400 ;
        RECT 1154.690 0.350 1157.270 1.400 ;
        RECT 1158.370 0.350 1160.950 1.400 ;
        RECT 1162.050 0.350 1164.630 1.400 ;
        RECT 1165.730 0.350 1168.310 1.400 ;
        RECT 1169.410 0.350 1171.990 1.400 ;
        RECT 1173.090 0.350 1175.670 1.400 ;
        RECT 1176.770 0.350 1179.350 1.400 ;
        RECT 1180.450 0.350 1183.030 1.400 ;
        RECT 1184.130 0.350 1194.990 1.400 ;
        RECT 1196.090 0.350 1198.670 1.400 ;
        RECT 1199.770 0.350 1202.350 1.400 ;
        RECT 1203.450 0.350 1206.030 1.400 ;
        RECT 1207.130 0.350 1209.710 1.400 ;
        RECT 1210.810 0.350 1213.390 1.400 ;
        RECT 1214.490 0.350 1217.070 1.400 ;
        RECT 1218.170 0.350 1220.750 1.400 ;
        RECT 1221.850 0.350 1224.430 1.400 ;
        RECT 1225.530 0.350 1228.110 1.400 ;
        RECT 1229.210 0.350 1231.790 1.400 ;
        RECT 1232.890 0.350 1235.470 1.400 ;
        RECT 1236.570 0.350 1239.150 1.400 ;
        RECT 1240.250 0.350 1242.830 1.400 ;
        RECT 1243.930 0.350 1246.510 1.400 ;
        RECT 1247.610 0.350 1250.190 1.400 ;
        RECT 1251.290 0.350 1253.870 1.400 ;
        RECT 1254.970 0.350 1257.550 1.400 ;
        RECT 1258.650 0.350 1261.230 1.400 ;
        RECT 1262.330 0.350 1264.910 1.400 ;
        RECT 1266.010 0.350 1268.590 1.400 ;
        RECT 1269.690 0.350 1272.270 1.400 ;
        RECT 1273.370 0.350 1275.950 1.400 ;
        RECT 1277.050 0.350 1279.630 1.400 ;
        RECT 1280.730 0.350 1283.310 1.400 ;
        RECT 1284.410 0.350 1286.990 1.400 ;
        RECT 1288.090 0.350 1290.670 1.400 ;
        RECT 1291.770 0.350 1294.350 1.400 ;
        RECT 1295.450 0.350 1298.030 1.400 ;
        RECT 1299.130 0.350 1301.710 1.400 ;
        RECT 1302.810 0.350 1305.390 1.400 ;
        RECT 1306.490 0.350 1309.070 1.400 ;
        RECT 1310.170 0.350 1312.750 1.400 ;
        RECT 1313.850 0.350 1316.430 1.400 ;
        RECT 1317.530 0.350 1320.110 1.400 ;
        RECT 1321.210 0.350 1323.790 1.400 ;
        RECT 1324.890 0.350 1327.470 1.400 ;
        RECT 1328.570 0.350 1331.150 1.400 ;
        RECT 1332.250 0.350 1334.830 1.400 ;
        RECT 1335.930 0.350 1338.510 1.400 ;
        RECT 1339.610 0.350 1342.190 1.400 ;
        RECT 1343.290 0.350 1345.870 1.400 ;
        RECT 1346.970 0.350 1349.550 1.400 ;
        RECT 1350.650 0.350 1353.230 1.400 ;
  END
END tt_mux
END LIBRARY

