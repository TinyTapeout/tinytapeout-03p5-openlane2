VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_apu_pulse
  CLASS BLOCK ;
  FOREIGN tt_um_apu_pulse ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 106.950 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 85.500 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 85.500 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 85.500 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 106.950 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 89.550 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 82.100 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 85.500 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 85.500 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 11.380 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 61.950 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 85.500 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 84.820 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 19.540 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 21.580 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 106.950 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 3.900 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 106.580 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 87.540 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 89.580 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 106.950 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 85.500 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 63.060 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 86.180 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 89.580 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 83.460 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 106.950 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 84.820 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 15.460 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 85.500 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 106.950 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 106.950 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 86.550 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 106.950 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 61.950 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 28.380 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 106.950 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 35.180 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 88.900 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 107.260 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 20.220 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 86.860 66.850 108.800 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.325 5.200 25.925 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.535 5.200 65.135 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.745 5.200 104.345 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.955 5.200 143.555 103.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.930 5.200 45.530 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.140 5.200 84.740 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.350 5.200 123.950 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.560 5.200 163.160 103.600 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 162.380 103.445 ;
      LAYER met1 ;
        RECT 0.070 1.400 167.830 108.760 ;
      LAYER met2 ;
        RECT 0.090 1.370 167.800 108.790 ;
      LAYER met3 ;
        RECT 0.065 2.215 167.170 107.265 ;
      LAYER met4 ;
        RECT 0.295 83.060 7.270 108.450 ;
        RECT 8.370 89.180 10.950 108.450 ;
        RECT 12.050 89.180 14.630 108.450 ;
        RECT 8.370 85.780 14.630 89.180 ;
        RECT 15.730 85.780 18.310 108.450 ;
        RECT 8.370 83.060 18.310 85.780 ;
        RECT 0.295 62.660 18.310 83.060 ;
        RECT 19.410 85.100 21.990 108.450 ;
        RECT 23.090 106.550 25.670 108.450 ;
        RECT 26.770 106.550 29.350 108.450 ;
        RECT 23.090 104.000 29.350 106.550 ;
        RECT 23.090 85.100 23.925 104.000 ;
        RECT 19.410 62.660 23.925 85.100 ;
        RECT 0.295 4.800 23.925 62.660 ;
        RECT 26.325 89.180 29.350 104.000 ;
        RECT 30.450 89.180 33.030 108.450 ;
        RECT 26.325 87.140 33.030 89.180 ;
        RECT 34.130 106.550 36.710 108.450 ;
        RECT 37.810 106.550 40.390 108.450 ;
        RECT 34.130 87.140 40.390 106.550 ;
        RECT 26.325 86.150 40.390 87.140 ;
        RECT 41.490 106.550 44.070 108.450 ;
        RECT 45.170 106.550 47.750 108.450 ;
        RECT 48.850 106.550 51.430 108.450 ;
        RECT 41.490 104.000 51.430 106.550 ;
        RECT 41.490 86.150 43.530 104.000 ;
        RECT 26.325 4.800 43.530 86.150 ;
        RECT 45.930 85.100 51.430 104.000 ;
        RECT 52.530 85.100 55.110 108.450 ;
        RECT 45.930 15.060 55.110 85.100 ;
        RECT 56.210 84.420 58.790 108.450 ;
        RECT 59.890 106.550 62.470 108.450 ;
        RECT 63.570 106.550 66.150 108.450 ;
        RECT 59.890 104.000 66.150 106.550 ;
        RECT 59.890 84.420 63.135 104.000 ;
        RECT 56.210 15.060 63.135 84.420 ;
        RECT 45.930 4.800 63.135 15.060 ;
        RECT 65.535 86.460 66.150 104.000 ;
        RECT 67.250 86.460 69.830 108.450 ;
        RECT 65.535 19.820 69.830 86.460 ;
        RECT 70.930 106.860 73.510 108.450 ;
        RECT 74.610 106.860 77.190 108.450 ;
        RECT 70.930 88.500 77.190 106.860 ;
        RECT 78.290 88.500 80.870 108.450 ;
        RECT 70.930 34.780 80.870 88.500 ;
        RECT 81.970 106.550 84.550 108.450 ;
        RECT 85.650 106.550 88.230 108.450 ;
        RECT 81.970 104.000 88.230 106.550 ;
        RECT 81.970 34.780 82.740 104.000 ;
        RECT 70.930 19.820 82.740 34.780 ;
        RECT 65.535 4.800 82.740 19.820 ;
        RECT 85.140 27.980 88.230 104.000 ;
        RECT 89.330 61.550 91.910 108.450 ;
        RECT 93.010 106.180 95.590 108.450 ;
        RECT 96.690 106.180 99.270 108.450 ;
        RECT 93.010 61.550 99.270 106.180 ;
        RECT 89.330 27.980 99.270 61.550 ;
        RECT 85.140 4.800 99.270 27.980 ;
        RECT 0.295 3.500 99.270 4.800 ;
        RECT 100.370 106.550 102.950 108.450 ;
        RECT 104.050 106.550 106.630 108.450 ;
        RECT 100.370 104.000 106.630 106.550 ;
        RECT 100.370 4.800 102.345 104.000 ;
        RECT 104.745 21.180 106.630 104.000 ;
        RECT 107.730 21.180 110.310 108.450 ;
        RECT 104.745 19.140 110.310 21.180 ;
        RECT 111.410 84.420 113.990 108.450 ;
        RECT 115.090 85.100 117.670 108.450 ;
        RECT 118.770 85.100 121.350 108.450 ;
        RECT 122.450 104.000 125.030 108.450 ;
        RECT 115.090 84.420 121.350 85.100 ;
        RECT 111.410 61.550 121.350 84.420 ;
        RECT 111.410 19.140 121.950 61.550 ;
        RECT 104.745 4.800 121.950 19.140 ;
        RECT 124.350 10.980 125.030 104.000 ;
        RECT 126.130 85.100 128.710 108.450 ;
        RECT 129.810 85.100 132.390 108.450 ;
        RECT 133.490 85.100 136.070 108.450 ;
        RECT 126.130 81.700 136.070 85.100 ;
        RECT 137.170 89.150 139.750 108.450 ;
        RECT 140.850 106.550 143.430 108.450 ;
        RECT 144.530 106.550 147.110 108.450 ;
        RECT 140.850 104.000 147.110 106.550 ;
        RECT 140.850 89.150 141.555 104.000 ;
        RECT 137.170 81.700 141.555 89.150 ;
        RECT 126.130 10.980 141.555 81.700 ;
        RECT 124.350 4.800 141.555 10.980 ;
        RECT 143.955 85.100 147.110 104.000 ;
        RECT 148.210 85.100 150.790 108.450 ;
        RECT 151.890 85.100 154.470 108.450 ;
        RECT 155.570 106.550 158.150 108.450 ;
        RECT 159.250 107.400 161.830 108.450 ;
        RECT 162.930 107.400 167.145 108.450 ;
        RECT 159.250 106.550 167.145 107.400 ;
        RECT 155.570 104.000 167.145 106.550 ;
        RECT 155.570 85.100 161.160 104.000 ;
        RECT 143.955 4.800 161.160 85.100 ;
        RECT 163.560 4.800 167.145 104.000 ;
        RECT 100.370 3.500 167.145 4.800 ;
        RECT 0.295 2.895 167.145 3.500 ;
  END
END tt_um_apu_pulse
END LIBRARY

