VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_ctrl
  CLASS BLOCK ;
  FOREIGN tt_ctrl ;
  ORIGIN 0.000 0.000 ;
  SIZE 185.840 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.610 2.480 25.210 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.710 2.480 90.310 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.810 2.480 155.410 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.310 2.480 21.910 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.410 2.480 87.010 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.510 2.480 152.110 109.040 ;
    END
  END VPWR
  PIN ctrl_ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 26.990 0.000 27.290 1.000 ;
    END
  END ctrl_ena
  PIN ctrl_sel_inc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 25.150 0.000 25.450 1.000 ;
    END
  END ctrl_sel_inc
  PIN ctrl_sel_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 23.310 0.000 23.610 1.000 ;
    END
  END ctrl_sel_rst_n
  PIN k_one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 19.630 0.000 19.930 1.000 ;
    END
  END k_one
  PIN k_zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 0.000 21.770 1.000 ;
    END
  END k_zero
  PIN pad_ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 164.990 0.000 165.290 1.000 ;
    END
  END pad_ui_in[0]
  PIN pad_ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 166.830 0.000 167.130 1.000 ;
    END
  END pad_ui_in[1]
  PIN pad_ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 180.630 110.520 180.930 111.520 ;
    END
  END pad_ui_in[2]
  PIN pad_ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 178.790 110.520 179.090 111.520 ;
    END
  END pad_ui_in[3]
  PIN pad_ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 176.950 110.520 177.250 111.520 ;
    END
  END pad_ui_in[4]
  PIN pad_ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 175.110 110.520 175.410 111.520 ;
    END
  END pad_ui_in[5]
  PIN pad_ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 173.270 110.520 173.570 111.520 ;
    END
  END pad_ui_in[6]
  PIN pad_ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 171.430 110.520 171.730 111.520 ;
    END
  END pad_ui_in[7]
  PIN pad_ui_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 169.590 110.520 169.890 111.520 ;
    END
  END pad_ui_in[8]
  PIN pad_ui_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 167.750 110.520 168.050 111.520 ;
    END
  END pad_ui_in[9]
  PIN pad_uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 30.670 110.520 30.970 111.520 ;
    END
  END pad_uio_in[0]
  PIN pad_uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 25.150 110.520 25.450 111.520 ;
    END
  END pad_uio_in[1]
  PIN pad_uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 19.630 110.520 19.930 111.520 ;
    END
  END pad_uio_in[2]
  PIN pad_uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 14.110 110.520 14.410 111.520 ;
    END
  END pad_uio_in[3]
  PIN pad_uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 8.590 110.520 8.890 111.520 ;
    END
  END pad_uio_in[4]
  PIN pad_uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 3.070 110.520 3.370 111.520 ;
    END
  END pad_uio_in[5]
  PIN pad_uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 8.590 0.000 8.890 1.000 ;
    END
  END pad_uio_in[6]
  PIN pad_uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 14.110 0.000 14.410 1.000 ;
    END
  END pad_uio_in[7]
  PIN pad_uio_oe_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 110.520 151.490 111.520 ;
    END
  END pad_uio_oe_n[0]
  PIN pad_uio_oe_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 28.830 110.520 29.130 111.520 ;
    END
  END pad_uio_oe_n[1]
  PIN pad_uio_oe_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 23.310 110.520 23.610 111.520 ;
    END
  END pad_uio_oe_n[2]
  PIN pad_uio_oe_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 17.790 110.520 18.090 111.520 ;
    END
  END pad_uio_oe_n[3]
  PIN pad_uio_oe_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 12.270 110.520 12.570 111.520 ;
    END
  END pad_uio_oe_n[4]
  PIN pad_uio_oe_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 6.750 110.520 7.050 111.520 ;
    END
  END pad_uio_oe_n[5]
  PIN pad_uio_oe_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 12.270 0.000 12.570 1.000 ;
    END
  END pad_uio_oe_n[6]
  PIN pad_uio_oe_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 17.790 0.000 18.090 1.000 ;
    END
  END pad_uio_oe_n[7]
  PIN pad_uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END pad_uio_out[0]
  PIN pad_uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END pad_uio_out[1]
  PIN pad_uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END pad_uio_out[2]
  PIN pad_uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 15.950 110.520 16.250 111.520 ;
    END
  END pad_uio_out[3]
  PIN pad_uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 10.430 110.520 10.730 111.520 ;
    END
  END pad_uio_out[4]
  PIN pad_uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 4.910 110.520 5.210 111.520 ;
    END
  END pad_uio_out[5]
  PIN pad_uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 10.430 0.000 10.730 1.000 ;
    END
  END pad_uio_out[6]
  PIN pad_uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 15.950 0.000 16.250 1.000 ;
    END
  END pad_uio_out[7]
  PIN pad_uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 165.910 110.520 166.210 111.520 ;
    END
  END pad_uo_out[0]
  PIN pad_uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 164.070 110.520 164.370 111.520 ;
    END
  END pad_uo_out[1]
  PIN pad_uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 162.230 110.520 162.530 111.520 ;
    END
  END pad_uo_out[2]
  PIN pad_uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 160.390 110.520 160.690 111.520 ;
    END
  END pad_uo_out[3]
  PIN pad_uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 158.550 110.520 158.850 111.520 ;
    END
  END pad_uo_out[4]
  PIN pad_uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 156.710 110.520 157.010 111.520 ;
    END
  END pad_uo_out[5]
  PIN pad_uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 110.520 155.170 111.520 ;
    END
  END pad_uo_out[6]
  PIN pad_uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 153.030 110.520 153.330 111.520 ;
    END
  END pad_uo_out[7]
  PIN spine_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 0.000 146.890 111.520 ;
    END
  END spine_iw[0]
  PIN spine_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 0.000 128.490 111.520 ;
    END
  END spine_iw[10]
  PIN spine_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 0.000 126.650 111.520 ;
    END
  END spine_iw[11]
  PIN spine_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 0.000 124.810 111.520 ;
    END
  END spine_iw[12]
  PIN spine_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 0.000 122.970 111.520 ;
    END
  END spine_iw[13]
  PIN spine_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 120.830 0.000 121.130 111.520 ;
    END
  END spine_iw[14]
  PIN spine_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 0.000 119.290 111.520 ;
    END
  END spine_iw[15]
  PIN spine_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 0.000 117.450 111.520 ;
    END
  END spine_iw[16]
  PIN spine_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 115.310 0.000 115.610 111.520 ;
    END
  END spine_iw[17]
  PIN spine_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 0.000 113.770 111.520 ;
    END
  END spine_iw[18]
  PIN spine_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 0.000 111.930 111.520 ;
    END
  END spine_iw[19]
  PIN spine_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 144.750 0.000 145.050 111.520 ;
    END
  END spine_iw[1]
  PIN spine_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 109.790 0.000 110.090 111.520 ;
    END
  END spine_iw[20]
  PIN spine_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 0.000 108.250 111.520 ;
    END
  END spine_iw[21]
  PIN spine_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 0.000 106.410 111.520 ;
    END
  END spine_iw[22]
  PIN spine_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 104.270 0.000 104.570 111.520 ;
    END
  END spine_iw[23]
  PIN spine_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 102.430 0.000 102.730 111.520 ;
    END
  END spine_iw[24]
  PIN spine_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 0.000 100.890 111.520 ;
    END
  END spine_iw[25]
  PIN spine_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 98.750 0.000 99.050 111.520 ;
    END
  END spine_iw[26]
  PIN spine_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 96.910 0.000 97.210 111.520 ;
    END
  END spine_iw[27]
  PIN spine_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 0.000 95.370 111.520 ;
    END
  END spine_iw[28]
  PIN spine_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 93.230 0.000 93.530 111.520 ;
    END
  END spine_iw[29]
  PIN spine_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 142.910 0.000 143.210 111.520 ;
    END
  END spine_iw[2]
  PIN spine_iw[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 0.000 91.690 111.520 ;
    END
  END spine_iw[30]
  PIN spine_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 0.000 141.370 111.520 ;
    END
  END spine_iw[3]
  PIN spine_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 139.230 0.000 139.530 111.520 ;
    END
  END spine_iw[4]
  PIN spine_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 137.390 0.000 137.690 111.520 ;
    END
  END spine_iw[5]
  PIN spine_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 0.000 135.850 111.520 ;
    END
  END spine_iw[6]
  PIN spine_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 133.710 0.000 134.010 111.520 ;
    END
  END spine_iw[7]
  PIN spine_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 131.870 0.000 132.170 111.520 ;
    END
  END spine_iw[8]
  PIN spine_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 0.000 130.330 111.520 ;
    END
  END spine_iw[9]
  PIN spine_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 0.000 84.330 111.520 ;
    END
  END spine_ow[0]
  PIN spine_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 65.630 0.000 65.930 111.520 ;
    END
  END spine_ow[10]
  PIN spine_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 0.000 64.090 111.520 ;
    END
  END spine_ow[11]
  PIN spine_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 0.000 62.250 111.520 ;
    END
  END spine_ow[12]
  PIN spine_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 60.110 0.000 60.410 111.520 ;
    END
  END spine_ow[13]
  PIN spine_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 58.270 0.000 58.570 111.520 ;
    END
  END spine_ow[14]
  PIN spine_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 56.430 0.000 56.730 111.520 ;
    END
  END spine_ow[15]
  PIN spine_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 54.590 0.000 54.890 111.520 ;
    END
  END spine_ow[16]
  PIN spine_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 52.750 0.000 53.050 111.520 ;
    END
  END spine_ow[17]
  PIN spine_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 50.910 0.000 51.210 111.520 ;
    END
  END spine_ow[18]
  PIN spine_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 49.070 0.000 49.370 111.520 ;
    END
  END spine_ow[19]
  PIN spine_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 82.190 0.000 82.490 111.520 ;
    END
  END spine_ow[1]
  PIN spine_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 47.230 0.000 47.530 111.520 ;
    END
  END spine_ow[20]
  PIN spine_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 45.390 0.000 45.690 111.520 ;
    END
  END spine_ow[21]
  PIN spine_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 43.550 0.000 43.850 111.520 ;
    END
  END spine_ow[22]
  PIN spine_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 41.710 0.000 42.010 111.520 ;
    END
  END spine_ow[23]
  PIN spine_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 39.870 0.000 40.170 111.520 ;
    END
  END spine_ow[24]
  PIN spine_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.030 0.000 38.330 111.520 ;
    END
  END spine_ow[25]
  PIN spine_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 0.000 80.650 111.520 ;
    END
  END spine_ow[2]
  PIN spine_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 0.000 78.810 111.520 ;
    END
  END spine_ow[3]
  PIN spine_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 76.670 0.000 76.970 111.520 ;
    END
  END spine_ow[4]
  PIN spine_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 0.000 75.130 111.520 ;
    END
  END spine_ow[5]
  PIN spine_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 0.000 73.290 111.520 ;
    END
  END spine_ow[6]
  PIN spine_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 71.150 0.000 71.450 111.520 ;
    END
  END spine_ow[7]
  PIN spine_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 0.000 69.610 111.520 ;
    END
  END spine_ow[8]
  PIN spine_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 0.000 67.770 111.520 ;
    END
  END spine_ow[9]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 183.270 108.990 ;
        RECT 2.570 101.945 183.270 104.775 ;
        RECT 2.570 96.505 183.270 99.335 ;
        RECT 2.570 91.065 183.270 93.895 ;
        RECT 2.570 85.625 183.270 88.455 ;
        RECT 2.570 80.185 183.270 83.015 ;
        RECT 2.570 74.745 183.270 77.575 ;
        RECT 2.570 69.305 183.270 72.135 ;
        RECT 2.570 63.865 183.270 66.695 ;
        RECT 2.570 58.425 183.270 61.255 ;
        RECT 2.570 52.985 183.270 55.815 ;
        RECT 2.570 47.545 183.270 50.375 ;
        RECT 2.570 42.105 183.270 44.935 ;
        RECT 2.570 36.665 183.270 39.495 ;
        RECT 2.570 31.225 183.270 34.055 ;
        RECT 2.570 25.785 183.270 28.615 ;
        RECT 2.570 20.345 183.270 23.175 ;
        RECT 2.570 14.905 183.270 17.735 ;
        RECT 2.570 9.465 183.270 12.295 ;
        RECT 2.570 4.025 183.270 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 183.080 108.885 ;
      LAYER met1 ;
        RECT 2.760 2.480 183.080 109.040 ;
      LAYER met2 ;
        RECT 5.150 1.515 174.250 110.005 ;
      LAYER met3 ;
        RECT 3.030 1.535 180.970 109.985 ;
      LAYER met4 ;
        RECT 3.770 110.120 4.510 111.170 ;
        RECT 5.610 110.120 6.350 111.170 ;
        RECT 7.450 110.120 8.190 111.170 ;
        RECT 9.290 110.120 10.030 111.170 ;
        RECT 11.130 110.120 11.870 111.170 ;
        RECT 12.970 110.120 13.710 111.170 ;
        RECT 14.810 110.120 15.550 111.170 ;
        RECT 16.650 110.120 17.390 111.170 ;
        RECT 18.490 110.120 19.230 111.170 ;
        RECT 20.330 110.120 21.070 111.170 ;
        RECT 22.170 110.120 22.910 111.170 ;
        RECT 24.010 110.120 24.750 111.170 ;
        RECT 25.850 110.120 26.590 111.170 ;
        RECT 27.690 110.120 28.430 111.170 ;
        RECT 29.530 110.120 30.270 111.170 ;
        RECT 31.370 110.120 32.110 111.170 ;
        RECT 33.210 110.120 37.630 111.170 ;
        RECT 3.055 109.440 37.630 110.120 ;
        RECT 3.055 2.080 19.910 109.440 ;
        RECT 22.310 2.080 23.210 109.440 ;
        RECT 25.610 2.080 37.630 109.440 ;
        RECT 3.055 1.400 37.630 2.080 ;
        RECT 3.055 1.000 8.190 1.400 ;
        RECT 9.290 1.000 10.030 1.400 ;
        RECT 11.130 1.000 11.870 1.400 ;
        RECT 12.970 1.000 13.710 1.400 ;
        RECT 14.810 1.000 15.550 1.400 ;
        RECT 16.650 1.000 17.390 1.400 ;
        RECT 18.490 1.000 19.230 1.400 ;
        RECT 20.330 1.000 21.070 1.400 ;
        RECT 22.170 1.000 22.910 1.400 ;
        RECT 24.010 1.000 24.750 1.400 ;
        RECT 25.850 1.000 26.590 1.400 ;
        RECT 27.690 1.000 37.630 1.400 ;
        RECT 38.730 1.000 39.470 111.170 ;
        RECT 40.570 1.000 41.310 111.170 ;
        RECT 42.410 1.000 43.150 111.170 ;
        RECT 44.250 1.000 44.990 111.170 ;
        RECT 46.090 1.000 46.830 111.170 ;
        RECT 47.930 1.000 48.670 111.170 ;
        RECT 49.770 1.000 50.510 111.170 ;
        RECT 51.610 1.000 52.350 111.170 ;
        RECT 53.450 1.000 54.190 111.170 ;
        RECT 55.290 1.000 56.030 111.170 ;
        RECT 57.130 1.000 57.870 111.170 ;
        RECT 58.970 1.000 59.710 111.170 ;
        RECT 60.810 1.000 61.550 111.170 ;
        RECT 62.650 1.000 63.390 111.170 ;
        RECT 64.490 1.000 65.230 111.170 ;
        RECT 66.330 1.000 67.070 111.170 ;
        RECT 68.170 1.000 68.910 111.170 ;
        RECT 70.010 1.000 70.750 111.170 ;
        RECT 71.850 1.000 72.590 111.170 ;
        RECT 73.690 1.000 74.430 111.170 ;
        RECT 75.530 1.000 76.270 111.170 ;
        RECT 77.370 1.000 78.110 111.170 ;
        RECT 79.210 1.000 79.950 111.170 ;
        RECT 81.050 1.000 81.790 111.170 ;
        RECT 82.890 1.000 83.630 111.170 ;
        RECT 84.730 109.440 90.990 111.170 ;
        RECT 84.730 2.080 85.010 109.440 ;
        RECT 87.410 2.080 88.310 109.440 ;
        RECT 90.710 2.080 90.990 109.440 ;
        RECT 84.730 1.000 90.990 2.080 ;
        RECT 92.090 1.000 92.830 111.170 ;
        RECT 93.930 1.000 94.670 111.170 ;
        RECT 95.770 1.000 96.510 111.170 ;
        RECT 97.610 1.000 98.350 111.170 ;
        RECT 99.450 1.000 100.190 111.170 ;
        RECT 101.290 1.000 102.030 111.170 ;
        RECT 103.130 1.000 103.870 111.170 ;
        RECT 104.970 1.000 105.710 111.170 ;
        RECT 106.810 1.000 107.550 111.170 ;
        RECT 108.650 1.000 109.390 111.170 ;
        RECT 110.490 1.000 111.230 111.170 ;
        RECT 112.330 1.000 113.070 111.170 ;
        RECT 114.170 1.000 114.910 111.170 ;
        RECT 116.010 1.000 116.750 111.170 ;
        RECT 117.850 1.000 118.590 111.170 ;
        RECT 119.690 1.000 120.430 111.170 ;
        RECT 121.530 1.000 122.270 111.170 ;
        RECT 123.370 1.000 124.110 111.170 ;
        RECT 125.210 1.000 125.950 111.170 ;
        RECT 127.050 1.000 127.790 111.170 ;
        RECT 128.890 1.000 129.630 111.170 ;
        RECT 130.730 1.000 131.470 111.170 ;
        RECT 132.570 1.000 133.310 111.170 ;
        RECT 134.410 1.000 135.150 111.170 ;
        RECT 136.250 1.000 136.990 111.170 ;
        RECT 138.090 1.000 138.830 111.170 ;
        RECT 139.930 1.000 140.670 111.170 ;
        RECT 141.770 1.000 142.510 111.170 ;
        RECT 143.610 1.000 144.350 111.170 ;
        RECT 145.450 1.000 146.190 111.170 ;
        RECT 147.290 110.120 150.790 111.170 ;
        RECT 151.890 110.120 152.630 111.170 ;
        RECT 153.730 110.120 154.470 111.170 ;
        RECT 155.570 110.120 156.310 111.170 ;
        RECT 157.410 110.120 158.150 111.170 ;
        RECT 159.250 110.120 159.990 111.170 ;
        RECT 161.090 110.120 161.830 111.170 ;
        RECT 162.930 110.120 163.670 111.170 ;
        RECT 164.770 110.120 165.510 111.170 ;
        RECT 166.610 110.120 167.350 111.170 ;
        RECT 168.450 110.120 169.190 111.170 ;
        RECT 170.290 110.120 171.030 111.170 ;
        RECT 172.130 110.120 172.870 111.170 ;
        RECT 173.970 110.120 174.710 111.170 ;
        RECT 175.810 110.120 176.550 111.170 ;
        RECT 177.650 110.120 178.390 111.170 ;
        RECT 179.490 110.120 180.230 111.170 ;
        RECT 147.290 109.440 180.945 110.120 ;
        RECT 147.290 2.080 150.110 109.440 ;
        RECT 152.510 2.080 153.410 109.440 ;
        RECT 155.810 2.080 180.945 109.440 ;
        RECT 147.290 1.400 180.945 2.080 ;
        RECT 147.290 1.000 164.590 1.400 ;
        RECT 165.690 1.000 166.430 1.400 ;
        RECT 167.530 1.000 180.945 1.400 ;
  END
END tt_ctrl
END LIBRARY

