VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_ringosc_cnt
  CLASS BLOCK ;
  FOREIGN tt_um_ringosc_cnt ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 107.800 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.800 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 89.580 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 103.180 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.260 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 106.580 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.260 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 107.260 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 107.260 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.260 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.800 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 107.800 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 107.800 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.800 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.800 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 107.800 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.800 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.800 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 100.460 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 107.260 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 104.540 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 100.460 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 102.500 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 102.500 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 102.500 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 100.460 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 101.820 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 107.260 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 107.260 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 101.140 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 106.580 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 107.260 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 107.260 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 107.260 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 107.260 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 107.260 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 107.260 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 106.580 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 107.260 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 107.260 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 84.820 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 107.260 66.850 108.800 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.325 5.200 25.925 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.535 5.200 65.135 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.745 5.200 104.345 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.955 5.200 143.555 103.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.930 5.200 45.530 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.140 5.200 84.740 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.350 5.200 123.950 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.560 5.200 163.160 103.600 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 99.225 162.570 102.055 ;
        RECT 5.330 93.785 162.570 96.615 ;
        RECT 5.330 88.345 162.570 91.175 ;
        RECT 5.330 82.905 162.570 85.735 ;
        RECT 5.330 77.465 162.570 80.295 ;
        RECT 5.330 72.025 162.570 74.855 ;
        RECT 5.330 66.585 162.570 69.415 ;
        RECT 5.330 61.145 162.570 63.975 ;
        RECT 5.330 55.705 162.570 58.535 ;
        RECT 5.330 50.265 162.570 53.095 ;
        RECT 5.330 44.825 162.570 47.655 ;
        RECT 5.330 39.385 162.570 42.215 ;
        RECT 5.330 33.945 162.570 36.775 ;
        RECT 5.330 28.505 162.570 31.335 ;
        RECT 5.330 23.065 162.570 25.895 ;
        RECT 5.330 17.625 162.570 20.455 ;
        RECT 5.330 12.185 162.570 15.015 ;
        RECT 5.330 6.745 162.570 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 162.380 103.445 ;
      LAYER met1 ;
        RECT 5.520 5.200 163.160 107.060 ;
      LAYER met2 ;
        RECT 7.910 5.255 163.130 107.285 ;
      LAYER met3 ;
        RECT 7.630 5.275 163.150 107.265 ;
      LAYER met4 ;
        RECT 8.370 102.100 10.950 107.265 ;
        RECT 12.050 102.100 14.630 107.265 ;
        RECT 15.730 102.100 18.310 107.265 ;
        RECT 19.410 102.100 21.990 107.265 ;
        RECT 8.370 100.060 21.990 102.100 ;
        RECT 23.090 104.140 25.670 107.265 ;
        RECT 26.770 106.860 29.350 107.265 ;
        RECT 30.450 106.860 33.030 107.265 ;
        RECT 26.770 104.140 33.030 106.860 ;
        RECT 23.090 104.000 33.030 104.140 ;
        RECT 23.090 100.060 23.925 104.000 ;
        RECT 7.655 57.295 23.925 100.060 ;
        RECT 26.325 100.060 33.030 104.000 ;
        RECT 34.130 106.860 36.710 107.265 ;
        RECT 37.810 106.860 40.390 107.265 ;
        RECT 41.490 106.860 44.070 107.265 ;
        RECT 45.170 106.860 47.750 107.265 ;
        RECT 34.130 106.180 47.750 106.860 ;
        RECT 48.850 106.180 51.430 107.265 ;
        RECT 34.130 104.000 51.430 106.180 ;
        RECT 34.130 100.060 43.530 104.000 ;
        RECT 26.325 57.295 43.530 100.060 ;
        RECT 45.930 100.740 51.430 104.000 ;
        RECT 52.530 106.860 55.110 107.265 ;
        RECT 56.210 106.860 58.790 107.265 ;
        RECT 59.890 106.860 62.470 107.265 ;
        RECT 52.530 101.420 62.470 106.860 ;
        RECT 63.570 106.860 66.150 107.265 ;
        RECT 67.250 106.860 69.830 107.265 ;
        RECT 63.570 104.000 69.830 106.860 ;
        RECT 52.530 100.740 63.135 101.420 ;
        RECT 45.930 57.295 63.135 100.740 ;
        RECT 65.535 84.420 69.830 104.000 ;
        RECT 70.930 106.860 73.510 107.265 ;
        RECT 74.610 106.860 77.190 107.265 ;
        RECT 78.290 106.860 80.870 107.265 ;
        RECT 70.930 106.180 80.870 106.860 ;
        RECT 81.970 106.860 84.550 107.265 ;
        RECT 85.650 106.860 88.230 107.265 ;
        RECT 89.330 106.860 91.910 107.265 ;
        RECT 93.010 106.860 125.030 107.265 ;
        RECT 126.130 106.860 128.710 107.265 ;
        RECT 129.810 106.860 132.390 107.265 ;
        RECT 133.490 106.860 136.070 107.265 ;
        RECT 137.170 106.860 139.750 107.265 ;
        RECT 81.970 106.180 139.750 106.860 ;
        RECT 140.850 106.860 143.430 107.265 ;
        RECT 144.530 106.860 147.110 107.265 ;
        RECT 140.850 106.180 147.110 106.860 ;
        RECT 70.930 104.000 147.110 106.180 ;
        RECT 70.930 84.420 82.740 104.000 ;
        RECT 65.535 57.295 82.740 84.420 ;
        RECT 85.140 57.295 102.345 104.000 ;
        RECT 104.745 57.295 121.950 104.000 ;
        RECT 124.350 57.295 141.555 104.000 ;
        RECT 143.955 102.780 147.110 104.000 ;
        RECT 148.210 102.780 150.790 107.265 ;
        RECT 143.955 89.180 150.790 102.780 ;
        RECT 143.955 57.295 151.505 89.180 ;
  END
END tt_um_ringosc_cnt
END LIBRARY

